// ROMs Using Block RAM Resources.
// File: rams_sp_rom_1.v
//
module background_rom(clk, en, addr, dout);
input clk;
input en;
input [13:0] addr;
output dout;

logic data;

always_ff @(posedge clk) begin
    if (en)
        case(addr)
0: data <= 'd0; 1: data <= 'd0; 2: data <= 'd0; 3: data <= 'd0; 4: data <= 'd0; 5: data <= 'd0; 6: data <= 'd0; 7: data <= 'd0; 8: data <= 'd0; 9: data <= 'd0; 10: data <= 'd0; 11: data <= 'd0; 12: data <= 'd0; 13: data <= 'd0; 14: data <= 'd0; 15: data <= 'd0; 16: data <= 'd0; 17: data <= 'd0; 18: data <= 'd0; 19: data <= 'd0; 20: data <= 'd0; 21: data <= 'd0; 22: data <= 'd0; 23: data <= 'd0; 24: data <= 'd0; 25: data <= 'd0; 26: data <= 'd0; 27: data <= 'd0; 28: data <= 'd0; 29: data <= 'd0; 30: data <= 'd0; 31: data <= 'd0; 32: data <= 'd0; 33: data <= 'd0; 34: data <= 'd0; 35: data <= 'd0; 36: data <= 'd0; 37: data <= 'd0; 38: data <= 'd0; 39: data <= 'd0; 40: data <= 'd0; 41: data <= 'd0; 42: data <= 'd0; 43: data <= 'd0; 44: data <= 'd0; 45: data <= 'd0; 46: data <= 'd0; 47: data <= 'd0; 48: data <= 'd0; 49: data <= 'd0; 50: data <= 'd0; 51: data <= 'd0; 52: data <= 'd0; 53: data <= 'd0; 54: data <= 'd0; 55: data <= 'd0; 56: data <= 'd0; 57: data <= 'd0; 58: data <= 'd0; 59: data <= 'd0; 60: data <= 'd0; 61: data <= 'd0; 62: data <= 'd0; 63: data <= 'd0; 64: data <= 'd0; 65: data <= 'd0; 66: data <= 'd0; 67: data <= 'd0; 68: data <= 'd0; 69: data <= 'd0; 70: data <= 'd0; 71: data <= 'd0; 72: data <= 'd0; 73: data <= 'd0; 74: data <= 'd0; 75: data <= 'd0; 76: data <= 'd0; 77: data <= 'd0; 78: data <= 'd0; 79: data <= 'd0; 80: data <= 'd0; 81: data <= 'd0; 82: data <= 'd0; 83: data <= 'd0; 84: data <= 'd0; 85: data <= 'd0; 86: data <= 'd0; 87: data <= 'd0; 88: data <= 'd0; 89: data <= 'd0; 90: data <= 'd0; 91: data <= 'd0; 92: data <= 'd0; 93: data <= 'd0; 94: data <= 'd0; 95: data <= 'd0; 96: data <= 'd0; 97: data <= 'd0; 98: data <= 'd0; 99: data <= 'd0; 100: data <= 'd0; 101: data <= 'd0; 102: data <= 'd0; 103: data <= 'd0; 104: data <= 'd0; 105: data <= 'd0; 106: data <= 'd0; 107: data <= 'd0; 108: data <= 'd0; 109: data <= 'd0; 110: data <= 'd0; 111: data <= 'd0; 112: data <= 'd0; 113: data <= 'd0; 114: data <= 'd0; 115: data <= 'd0; 116: data <= 'd0; 117: data <= 'd0; 118: data <= 'd0; 119: data <= 'd0; 120: data <= 'd0; 121: data <= 'd0; 122: data <= 'd0; 123: data <= 'd0; 124: data <= 'd0; 125: data <= 'd0; 126: data <= 'd0; 127: data <= 'd1; 128: data <= 'd0; 129: data <= 'd0; 130: data <= 'd0; 131: data <= 'd0; 132: data <= 'd0; 133: data <= 'd0; 134: data <= 'd0; 135: data <= 'd0; 136: data <= 'd0; 137: data <= 'd0; 138: data <= 'd0; 139: data <= 'd0; 140: data <= 'd0; 141: data <= 'd0; 142: data <= 'd0; 143: data <= 'd0; 144: data <= 'd0; 145: data <= 'd0; 146: data <= 'd0; 147: data <= 'd0; 148: data <= 'd0; 149: data <= 'd0; 150: data <= 'd0; 151: data <= 'd0; 152: data <= 'd0; 153: data <= 'd0; 154: data <= 'd0; 155: data <= 'd0; 156: data <= 'd0; 157: data <= 'd0; 158: data <= 'd0; 159: data <= 'd0; 160: data <= 'd0; 161: data <= 'd0; 162: data <= 'd0; 163: data <= 'd0; 164: data <= 'd0; 165: data <= 'd0; 166: data <= 'd0; 167: data <= 'd0; 168: data <= 'd0; 169: data <= 'd0; 170: data <= 'd0; 171: data <= 'd0; 172: data <= 'd0; 173: data <= 'd0; 174: data <= 'd0; 175: data <= 'd0; 176: data <= 'd0; 177: data <= 'd0; 178: data <= 'd0; 179: data <= 'd0; 180: data <= 'd0; 181: data <= 'd0; 182: data <= 'd0; 183: data <= 'd0; 184: data <= 'd0; 185: data <= 'd0; 186: data <= 'd0; 187: data <= 'd0; 188: data <= 'd0; 189: data <= 'd0; 190: data <= 'd0; 191: data <= 'd0; 192: data <= 'd0; 193: data <= 'd0; 194: data <= 'd0; 195: data <= 'd0; 196: data <= 'd0; 197: data <= 'd0; 198: data <= 'd0; 199: data <= 'd0; 200: data <= 'd0; 201: data <= 'd0; 202: data <= 'd0; 203: data <= 'd0; 204: data <= 'd0; 205: data <= 'd0; 206: data <= 'd0; 207: data <= 'd0; 208: data <= 'd0; 209: data <= 'd0; 210: data <= 'd0; 211: data <= 'd0; 212: data <= 'd0; 213: data <= 'd0; 214: data <= 'd0; 215: data <= 'd0; 216: data <= 'd0; 217: data <= 'd0; 218: data <= 'd0; 219: data <= 'd0; 220: data <= 'd0; 221: data <= 'd0; 222: data <= 'd0; 223: data <= 'd0; 224: data <= 'd0; 225: data <= 'd0; 226: data <= 'd0; 227: data <= 'd0; 228: data <= 'd0; 229: data <= 'd0; 230: data <= 'd0; 231: data <= 'd0; 232: data <= 'd0; 233: data <= 'd0; 234: data <= 'd0; 235: data <= 'd0; 236: data <= 'd0; 237: data <= 'd0; 238: data <= 'd0; 239: data <= 'd0; 240: data <= 'd0; 241: data <= 'd0; 242: data <= 'd0; 243: data <= 'd0; 244: data <= 'd0; 245: data <= 'd0; 246: data <= 'd0; 247: data <= 'd0; 248: data <= 'd0; 249: data <= 'd0; 250: data <= 'd0; 251: data <= 'd0; 252: data <= 'd0; 253: data <= 'd0; 254: data <= 'd0; 255: data <= 'd1; 256: data <= 'd0; 257: data <= 'd0; 258: data <= 'd0; 259: data <= 'd0; 260: data <= 'd0; 261: data <= 'd0; 262: data <= 'd0; 263: data <= 'd0; 264: data <= 'd0; 265: data <= 'd0; 266: data <= 'd0; 267: data <= 'd0; 268: data <= 'd0; 269: data <= 'd0; 270: data <= 'd0; 271: data <= 'd0; 272: data <= 'd0; 273: data <= 'd0; 274: data <= 'd0; 275: data <= 'd0; 276: data <= 'd0; 277: data <= 'd0; 278: data <= 'd0; 279: data <= 'd0; 280: data <= 'd0; 281: data <= 'd0; 282: data <= 'd0; 283: data <= 'd0; 284: data <= 'd0; 285: data <= 'd0; 286: data <= 'd0; 287: data <= 'd0; 288: data <= 'd0; 289: data <= 'd0; 290: data <= 'd0; 291: data <= 'd0; 292: data <= 'd0; 293: data <= 'd0; 294: data <= 'd0; 295: data <= 'd0; 296: data <= 'd0; 297: data <= 'd0; 298: data <= 'd0; 299: data <= 'd0; 300: data <= 'd0; 301: data <= 'd0; 302: data <= 'd0; 303: data <= 'd0; 304: data <= 'd0; 305: data <= 'd0; 306: data <= 'd0; 307: data <= 'd0; 308: data <= 'd0; 309: data <= 'd0; 310: data <= 'd0; 311: data <= 'd0; 312: data <= 'd0; 313: data <= 'd0; 314: data <= 'd0; 315: data <= 'd0; 316: data <= 'd0; 317: data <= 'd0; 318: data <= 'd0; 319: data <= 'd0; 320: data <= 'd0; 321: data <= 'd0; 322: data <= 'd0; 323: data <= 'd0; 324: data <= 'd0; 325: data <= 'd0; 326: data <= 'd0; 327: data <= 'd0; 328: data <= 'd0; 329: data <= 'd0; 330: data <= 'd0; 331: data <= 'd0; 332: data <= 'd0; 333: data <= 'd0; 334: data <= 'd0; 335: data <= 'd0; 336: data <= 'd0; 337: data <= 'd0; 338: data <= 'd0; 339: data <= 'd0; 340: data <= 'd0; 341: data <= 'd0; 342: data <= 'd0; 343: data <= 'd0; 344: data <= 'd0; 345: data <= 'd0; 346: data <= 'd0; 347: data <= 'd0; 348: data <= 'd0; 349: data <= 'd0; 350: data <= 'd0; 351: data <= 'd0; 352: data <= 'd0; 353: data <= 'd0; 354: data <= 'd0; 355: data <= 'd0; 356: data <= 'd0; 357: data <= 'd0; 358: data <= 'd0; 359: data <= 'd0; 360: data <= 'd0; 361: data <= 'd0; 362: data <= 'd0; 363: data <= 'd0; 364: data <= 'd0; 365: data <= 'd0; 366: data <= 'd0; 367: data <= 'd0; 368: data <= 'd0; 369: data <= 'd0; 370: data <= 'd0; 371: data <= 'd0; 372: data <= 'd0; 373: data <= 'd0; 374: data <= 'd0; 375: data <= 'd0; 376: data <= 'd0; 377: data <= 'd0; 378: data <= 'd0; 379: data <= 'd0; 380: data <= 'd0; 381: data <= 'd0; 382: data <= 'd0; 383: data <= 'd1; 384: data <= 'd0; 385: data <= 'd0; 386: data <= 'd0; 387: data <= 'd0; 388: data <= 'd0; 389: data <= 'd0; 390: data <= 'd0; 391: data <= 'd0; 392: data <= 'd0; 393: data <= 'd0; 394: data <= 'd0; 395: data <= 'd0; 396: data <= 'd0; 397: data <= 'd0; 398: data <= 'd0; 399: data <= 'd0; 400: data <= 'd0; 401: data <= 'd0; 402: data <= 'd0; 403: data <= 'd0; 404: data <= 'd0; 405: data <= 'd0; 406: data <= 'd0; 407: data <= 'd0; 408: data <= 'd0; 409: data <= 'd1; 410: data <= 'd1; 411: data <= 'd0; 412: data <= 'd0; 413: data <= 'd0; 414: data <= 'd0; 415: data <= 'd0; 416: data <= 'd0; 417: data <= 'd0; 418: data <= 'd0; 419: data <= 'd0; 420: data <= 'd0; 421: data <= 'd0; 422: data <= 'd0; 423: data <= 'd0; 424: data <= 'd0; 425: data <= 'd0; 426: data <= 'd0; 427: data <= 'd0; 428: data <= 'd0; 429: data <= 'd0; 430: data <= 'd0; 431: data <= 'd0; 432: data <= 'd0; 433: data <= 'd0; 434: data <= 'd0; 435: data <= 'd0; 436: data <= 'd0; 437: data <= 'd0; 438: data <= 'd0; 439: data <= 'd0; 440: data <= 'd0; 441: data <= 'd0; 442: data <= 'd0; 443: data <= 'd0; 444: data <= 'd0; 445: data <= 'd0; 446: data <= 'd0; 447: data <= 'd0; 448: data <= 'd0; 449: data <= 'd0; 450: data <= 'd0; 451: data <= 'd0; 452: data <= 'd0; 453: data <= 'd0; 454: data <= 'd0; 455: data <= 'd0; 456: data <= 'd0; 457: data <= 'd0; 458: data <= 'd0; 459: data <= 'd0; 460: data <= 'd0; 461: data <= 'd0; 462: data <= 'd0; 463: data <= 'd0; 464: data <= 'd0; 465: data <= 'd0; 466: data <= 'd0; 467: data <= 'd0; 468: data <= 'd0; 469: data <= 'd0; 470: data <= 'd0; 471: data <= 'd0; 472: data <= 'd0; 473: data <= 'd0; 474: data <= 'd0; 475: data <= 'd0; 476: data <= 'd0; 477: data <= 'd0; 478: data <= 'd0; 479: data <= 'd0; 480: data <= 'd0; 481: data <= 'd0; 482: data <= 'd0; 483: data <= 'd0; 484: data <= 'd0; 485: data <= 'd0; 486: data <= 'd0; 487: data <= 'd0; 488: data <= 'd0; 489: data <= 'd0; 490: data <= 'd0; 491: data <= 'd0; 492: data <= 'd0; 493: data <= 'd0; 494: data <= 'd0; 495: data <= 'd0; 496: data <= 'd0; 497: data <= 'd0; 498: data <= 'd0; 499: data <= 'd0; 500: data <= 'd0; 501: data <= 'd0; 502: data <= 'd0; 503: data <= 'd0; 504: data <= 'd0; 505: data <= 'd0; 506: data <= 'd0; 507: data <= 'd0; 508: data <= 'd0; 509: data <= 'd0; 510: data <= 'd1; 511: data <= 'd1; 512: data <= 'd0; 513: data <= 'd0; 514: data <= 'd0; 515: data <= 'd0; 516: data <= 'd0; 517: data <= 'd0; 518: data <= 'd0; 519: data <= 'd0; 520: data <= 'd0; 521: data <= 'd0; 522: data <= 'd0; 523: data <= 'd0; 524: data <= 'd0; 525: data <= 'd0; 526: data <= 'd0; 527: data <= 'd0; 528: data <= 'd0; 529: data <= 'd0; 530: data <= 'd0; 531: data <= 'd0; 532: data <= 'd0; 533: data <= 'd0; 534: data <= 'd0; 535: data <= 'd0; 536: data <= 'd1; 537: data <= 'd1; 538: data <= 'd1; 539: data <= 'd0; 540: data <= 'd0; 541: data <= 'd0; 542: data <= 'd0; 543: data <= 'd0; 544: data <= 'd0; 545: data <= 'd0; 546: data <= 'd0; 547: data <= 'd0; 548: data <= 'd0; 549: data <= 'd0; 550: data <= 'd0; 551: data <= 'd0; 552: data <= 'd0; 553: data <= 'd0; 554: data <= 'd0; 555: data <= 'd0; 556: data <= 'd0; 557: data <= 'd0; 558: data <= 'd0; 559: data <= 'd0; 560: data <= 'd0; 561: data <= 'd0; 562: data <= 'd0; 563: data <= 'd0; 564: data <= 'd0; 565: data <= 'd0; 566: data <= 'd0; 567: data <= 'd0; 568: data <= 'd0; 569: data <= 'd0; 570: data <= 'd0; 571: data <= 'd0; 572: data <= 'd0; 573: data <= 'd0; 574: data <= 'd0; 575: data <= 'd0; 576: data <= 'd0; 577: data <= 'd0; 578: data <= 'd0; 579: data <= 'd0; 580: data <= 'd0; 581: data <= 'd0; 582: data <= 'd0; 583: data <= 'd0; 584: data <= 'd0; 585: data <= 'd0; 586: data <= 'd0; 587: data <= 'd0; 588: data <= 'd0; 589: data <= 'd0; 590: data <= 'd0; 591: data <= 'd0; 592: data <= 'd0; 593: data <= 'd0; 594: data <= 'd0; 595: data <= 'd0; 596: data <= 'd0; 597: data <= 'd0; 598: data <= 'd0; 599: data <= 'd0; 600: data <= 'd0; 601: data <= 'd0; 602: data <= 'd0; 603: data <= 'd0; 604: data <= 'd0; 605: data <= 'd0; 606: data <= 'd0; 607: data <= 'd0; 608: data <= 'd0; 609: data <= 'd0; 610: data <= 'd0; 611: data <= 'd0; 612: data <= 'd0; 613: data <= 'd0; 614: data <= 'd0; 615: data <= 'd0; 616: data <= 'd0; 617: data <= 'd0; 618: data <= 'd0; 619: data <= 'd0; 620: data <= 'd0; 621: data <= 'd0; 622: data <= 'd0; 623: data <= 'd0; 624: data <= 'd0; 625: data <= 'd0; 626: data <= 'd0; 627: data <= 'd0; 628: data <= 'd0; 629: data <= 'd0; 630: data <= 'd0; 631: data <= 'd0; 632: data <= 'd0; 633: data <= 'd0; 634: data <= 'd0; 635: data <= 'd0; 636: data <= 'd0; 637: data <= 'd0; 638: data <= 'd1; 639: data <= 'd1; 640: data <= 'd0; 641: data <= 'd0; 642: data <= 'd0; 643: data <= 'd0; 644: data <= 'd0; 645: data <= 'd0; 646: data <= 'd0; 647: data <= 'd0; 648: data <= 'd0; 649: data <= 'd0; 650: data <= 'd0; 651: data <= 'd0; 652: data <= 'd0; 653: data <= 'd0; 654: data <= 'd0; 655: data <= 'd0; 656: data <= 'd0; 657: data <= 'd0; 658: data <= 'd0; 659: data <= 'd0; 660: data <= 'd0; 661: data <= 'd0; 662: data <= 'd0; 663: data <= 'd1; 664: data <= 'd1; 665: data <= 'd1; 666: data <= 'd0; 667: data <= 'd0; 668: data <= 'd0; 669: data <= 'd0; 670: data <= 'd0; 671: data <= 'd0; 672: data <= 'd0; 673: data <= 'd0; 674: data <= 'd0; 675: data <= 'd0; 676: data <= 'd0; 677: data <= 'd0; 678: data <= 'd0; 679: data <= 'd0; 680: data <= 'd0; 681: data <= 'd0; 682: data <= 'd0; 683: data <= 'd0; 684: data <= 'd0; 685: data <= 'd0; 686: data <= 'd0; 687: data <= 'd0; 688: data <= 'd0; 689: data <= 'd0; 690: data <= 'd0; 691: data <= 'd0; 692: data <= 'd0; 693: data <= 'd0; 694: data <= 'd0; 695: data <= 'd0; 696: data <= 'd0; 697: data <= 'd0; 698: data <= 'd0; 699: data <= 'd0; 700: data <= 'd0; 701: data <= 'd0; 702: data <= 'd0; 703: data <= 'd0; 704: data <= 'd0; 705: data <= 'd0; 706: data <= 'd0; 707: data <= 'd0; 708: data <= 'd0; 709: data <= 'd0; 710: data <= 'd0; 711: data <= 'd0; 712: data <= 'd0; 713: data <= 'd0; 714: data <= 'd0; 715: data <= 'd0; 716: data <= 'd0; 717: data <= 'd0; 718: data <= 'd0; 719: data <= 'd0; 720: data <= 'd0; 721: data <= 'd0; 722: data <= 'd0; 723: data <= 'd0; 724: data <= 'd0; 725: data <= 'd0; 726: data <= 'd0; 727: data <= 'd0; 728: data <= 'd0; 729: data <= 'd0; 730: data <= 'd0; 731: data <= 'd0; 732: data <= 'd0; 733: data <= 'd0; 734: data <= 'd0; 735: data <= 'd0; 736: data <= 'd0; 737: data <= 'd0; 738: data <= 'd0; 739: data <= 'd0; 740: data <= 'd0; 741: data <= 'd0; 742: data <= 'd0; 743: data <= 'd0; 744: data <= 'd0; 745: data <= 'd0; 746: data <= 'd0; 747: data <= 'd0; 748: data <= 'd0; 749: data <= 'd0; 750: data <= 'd0; 751: data <= 'd0; 752: data <= 'd0; 753: data <= 'd0; 754: data <= 'd0; 755: data <= 'd0; 756: data <= 'd0; 757: data <= 'd0; 758: data <= 'd0; 759: data <= 'd0; 760: data <= 'd0; 761: data <= 'd0; 762: data <= 'd0; 763: data <= 'd0; 764: data <= 'd0; 765: data <= 'd0; 766: data <= 'd1; 767: data <= 'd1; 768: data <= 'd0; 769: data <= 'd0; 770: data <= 'd0; 771: data <= 'd0; 772: data <= 'd0; 773: data <= 'd0; 774: data <= 'd0; 775: data <= 'd0; 776: data <= 'd0; 777: data <= 'd0; 778: data <= 'd0; 779: data <= 'd0; 780: data <= 'd0; 781: data <= 'd0; 782: data <= 'd0; 783: data <= 'd0; 784: data <= 'd0; 785: data <= 'd0; 786: data <= 'd0; 787: data <= 'd0; 788: data <= 'd0; 789: data <= 'd0; 790: data <= 'd0; 791: data <= 'd1; 792: data <= 'd1; 793: data <= 'd1; 794: data <= 'd0; 795: data <= 'd0; 796: data <= 'd0; 797: data <= 'd0; 798: data <= 'd0; 799: data <= 'd0; 800: data <= 'd0; 801: data <= 'd0; 802: data <= 'd0; 803: data <= 'd0; 804: data <= 'd0; 805: data <= 'd0; 806: data <= 'd0; 807: data <= 'd0; 808: data <= 'd0; 809: data <= 'd0; 810: data <= 'd0; 811: data <= 'd0; 812: data <= 'd0; 813: data <= 'd0; 814: data <= 'd0; 815: data <= 'd0; 816: data <= 'd0; 817: data <= 'd0; 818: data <= 'd0; 819: data <= 'd0; 820: data <= 'd0; 821: data <= 'd0; 822: data <= 'd0; 823: data <= 'd0; 824: data <= 'd0; 825: data <= 'd0; 826: data <= 'd0; 827: data <= 'd0; 828: data <= 'd0; 829: data <= 'd0; 830: data <= 'd0; 831: data <= 'd0; 832: data <= 'd0; 833: data <= 'd0; 834: data <= 'd0; 835: data <= 'd0; 836: data <= 'd0; 837: data <= 'd0; 838: data <= 'd0; 839: data <= 'd0; 840: data <= 'd0; 841: data <= 'd0; 842: data <= 'd0; 843: data <= 'd0; 844: data <= 'd0; 845: data <= 'd0; 846: data <= 'd0; 847: data <= 'd0; 848: data <= 'd0; 849: data <= 'd0; 850: data <= 'd0; 851: data <= 'd0; 852: data <= 'd0; 853: data <= 'd0; 854: data <= 'd0; 855: data <= 'd0; 856: data <= 'd0; 857: data <= 'd0; 858: data <= 'd0; 859: data <= 'd0; 860: data <= 'd0; 861: data <= 'd0; 862: data <= 'd0; 863: data <= 'd0; 864: data <= 'd0; 865: data <= 'd0; 866: data <= 'd0; 867: data <= 'd0; 868: data <= 'd0; 869: data <= 'd0; 870: data <= 'd0; 871: data <= 'd0; 872: data <= 'd0; 873: data <= 'd0; 874: data <= 'd0; 875: data <= 'd0; 876: data <= 'd0; 877: data <= 'd0; 878: data <= 'd0; 879: data <= 'd0; 880: data <= 'd0; 881: data <= 'd0; 882: data <= 'd0; 883: data <= 'd0; 884: data <= 'd0; 885: data <= 'd0; 886: data <= 'd0; 887: data <= 'd0; 888: data <= 'd0; 889: data <= 'd0; 890: data <= 'd0; 891: data <= 'd0; 892: data <= 'd0; 893: data <= 'd1; 894: data <= 'd1; 895: data <= 'd1; 896: data <= 'd0; 897: data <= 'd0; 898: data <= 'd0; 899: data <= 'd0; 900: data <= 'd0; 901: data <= 'd0; 902: data <= 'd0; 903: data <= 'd0; 904: data <= 'd0; 905: data <= 'd0; 906: data <= 'd0; 907: data <= 'd0; 908: data <= 'd0; 909: data <= 'd0; 910: data <= 'd0; 911: data <= 'd1; 912: data <= 'd1; 913: data <= 'd1; 914: data <= 'd0; 915: data <= 'd0; 916: data <= 'd0; 917: data <= 'd0; 918: data <= 'd0; 919: data <= 'd1; 920: data <= 'd1; 921: data <= 'd1; 922: data <= 'd0; 923: data <= 'd0; 924: data <= 'd0; 925: data <= 'd0; 926: data <= 'd0; 927: data <= 'd0; 928: data <= 'd0; 929: data <= 'd0; 930: data <= 'd0; 931: data <= 'd0; 932: data <= 'd0; 933: data <= 'd0; 934: data <= 'd0; 935: data <= 'd0; 936: data <= 'd0; 937: data <= 'd0; 938: data <= 'd0; 939: data <= 'd0; 940: data <= 'd0; 941: data <= 'd0; 942: data <= 'd0; 943: data <= 'd0; 944: data <= 'd0; 945: data <= 'd0; 946: data <= 'd0; 947: data <= 'd0; 948: data <= 'd0; 949: data <= 'd0; 950: data <= 'd0; 951: data <= 'd0; 952: data <= 'd0; 953: data <= 'd0; 954: data <= 'd0; 955: data <= 'd0; 956: data <= 'd0; 957: data <= 'd0; 958: data <= 'd0; 959: data <= 'd0; 960: data <= 'd0; 961: data <= 'd0; 962: data <= 'd0; 963: data <= 'd0; 964: data <= 'd0; 965: data <= 'd0; 966: data <= 'd0; 967: data <= 'd0; 968: data <= 'd0; 969: data <= 'd0; 970: data <= 'd0; 971: data <= 'd0; 972: data <= 'd0; 973: data <= 'd0; 974: data <= 'd0; 975: data <= 'd0; 976: data <= 'd0; 977: data <= 'd0; 978: data <= 'd0; 979: data <= 'd0; 980: data <= 'd0; 981: data <= 'd0; 982: data <= 'd0; 983: data <= 'd0; 984: data <= 'd0; 985: data <= 'd0; 986: data <= 'd0; 987: data <= 'd0; 988: data <= 'd0; 989: data <= 'd0; 990: data <= 'd0; 991: data <= 'd0; 992: data <= 'd0; 993: data <= 'd0; 994: data <= 'd0; 995: data <= 'd0; 996: data <= 'd0; 997: data <= 'd0; 998: data <= 'd0; 999: data <= 'd0; 1000: data <= 'd0; 1001: data <= 'd0; 1002: data <= 'd0; 1003: data <= 'd0; 1004: data <= 'd0; 1005: data <= 'd0; 1006: data <= 'd0; 1007: data <= 'd0; 1008: data <= 'd0; 1009: data <= 'd0; 1010: data <= 'd0; 1011: data <= 'd0; 1012: data <= 'd0; 1013: data <= 'd0; 1014: data <= 'd0; 1015: data <= 'd0; 1016: data <= 'd0; 1017: data <= 'd0; 1018: data <= 'd0; 1019: data <= 'd0; 1020: data <= 'd0; 1021: data <= 'd1; 1022: data <= 'd1; 1023: data <= 'd1; 1024: data <= 'd0; 1025: data <= 'd0; 1026: data <= 'd0; 1027: data <= 'd0; 1028: data <= 'd0; 1029: data <= 'd0; 1030: data <= 'd0; 1031: data <= 'd0; 1032: data <= 'd0; 1033: data <= 'd0; 1034: data <= 'd0; 1035: data <= 'd0; 1036: data <= 'd0; 1037: data <= 'd0; 1038: data <= 'd0; 1039: data <= 'd0; 1040: data <= 'd0; 1041: data <= 'd1; 1042: data <= 'd1; 1043: data <= 'd0; 1044: data <= 'd0; 1045: data <= 'd0; 1046: data <= 'd0; 1047: data <= 'd1; 1048: data <= 'd1; 1049: data <= 'd1; 1050: data <= 'd0; 1051: data <= 'd0; 1052: data <= 'd0; 1053: data <= 'd0; 1054: data <= 'd0; 1055: data <= 'd0; 1056: data <= 'd0; 1057: data <= 'd0; 1058: data <= 'd0; 1059: data <= 'd0; 1060: data <= 'd0; 1061: data <= 'd0; 1062: data <= 'd0; 1063: data <= 'd0; 1064: data <= 'd0; 1065: data <= 'd0; 1066: data <= 'd0; 1067: data <= 'd0; 1068: data <= 'd0; 1069: data <= 'd0; 1070: data <= 'd0; 1071: data <= 'd0; 1072: data <= 'd0; 1073: data <= 'd0; 1074: data <= 'd0; 1075: data <= 'd0; 1076: data <= 'd0; 1077: data <= 'd0; 1078: data <= 'd0; 1079: data <= 'd0; 1080: data <= 'd0; 1081: data <= 'd0; 1082: data <= 'd0; 1083: data <= 'd0; 1084: data <= 'd0; 1085: data <= 'd0; 1086: data <= 'd0; 1087: data <= 'd0; 1088: data <= 'd0; 1089: data <= 'd0; 1090: data <= 'd0; 1091: data <= 'd0; 1092: data <= 'd0; 1093: data <= 'd0; 1094: data <= 'd0; 1095: data <= 'd0; 1096: data <= 'd0; 1097: data <= 'd0; 1098: data <= 'd0; 1099: data <= 'd0; 1100: data <= 'd0; 1101: data <= 'd0; 1102: data <= 'd0; 1103: data <= 'd0; 1104: data <= 'd0; 1105: data <= 'd0; 1106: data <= 'd0; 1107: data <= 'd0; 1108: data <= 'd0; 1109: data <= 'd0; 1110: data <= 'd0; 1111: data <= 'd0; 1112: data <= 'd0; 1113: data <= 'd0; 1114: data <= 'd0; 1115: data <= 'd0; 1116: data <= 'd0; 1117: data <= 'd0; 1118: data <= 'd0; 1119: data <= 'd0; 1120: data <= 'd0; 1121: data <= 'd0; 1122: data <= 'd0; 1123: data <= 'd0; 1124: data <= 'd0; 1125: data <= 'd0; 1126: data <= 'd0; 1127: data <= 'd0; 1128: data <= 'd0; 1129: data <= 'd0; 1130: data <= 'd0; 1131: data <= 'd0; 1132: data <= 'd0; 1133: data <= 'd0; 1134: data <= 'd0; 1135: data <= 'd0; 1136: data <= 'd0; 1137: data <= 'd0; 1138: data <= 'd0; 1139: data <= 'd0; 1140: data <= 'd0; 1141: data <= 'd0; 1142: data <= 'd0; 1143: data <= 'd0; 1144: data <= 'd0; 1145: data <= 'd0; 1146: data <= 'd0; 1147: data <= 'd0; 1148: data <= 'd1; 1149: data <= 'd1; 1150: data <= 'd1; 1151: data <= 'd1; 1152: data <= 'd0; 1153: data <= 'd0; 1154: data <= 'd0; 1155: data <= 'd0; 1156: data <= 'd0; 1157: data <= 'd0; 1158: data <= 'd0; 1159: data <= 'd0; 1160: data <= 'd0; 1161: data <= 'd0; 1162: data <= 'd0; 1163: data <= 'd0; 1164: data <= 'd0; 1165: data <= 'd0; 1166: data <= 'd0; 1167: data <= 'd0; 1168: data <= 'd0; 1169: data <= 'd0; 1170: data <= 'd1; 1171: data <= 'd1; 1172: data <= 'd1; 1173: data <= 'd1; 1174: data <= 'd1; 1175: data <= 'd1; 1176: data <= 'd1; 1177: data <= 'd1; 1178: data <= 'd1; 1179: data <= 'd0; 1180: data <= 'd0; 1181: data <= 'd0; 1182: data <= 'd0; 1183: data <= 'd0; 1184: data <= 'd0; 1185: data <= 'd0; 1186: data <= 'd0; 1187: data <= 'd0; 1188: data <= 'd0; 1189: data <= 'd0; 1190: data <= 'd0; 1191: data <= 'd0; 1192: data <= 'd0; 1193: data <= 'd0; 1194: data <= 'd0; 1195: data <= 'd0; 1196: data <= 'd0; 1197: data <= 'd0; 1198: data <= 'd0; 1199: data <= 'd0; 1200: data <= 'd0; 1201: data <= 'd0; 1202: data <= 'd0; 1203: data <= 'd0; 1204: data <= 'd0; 1205: data <= 'd0; 1206: data <= 'd0; 1207: data <= 'd0; 1208: data <= 'd0; 1209: data <= 'd0; 1210: data <= 'd0; 1211: data <= 'd0; 1212: data <= 'd0; 1213: data <= 'd0; 1214: data <= 'd0; 1215: data <= 'd0; 1216: data <= 'd0; 1217: data <= 'd0; 1218: data <= 'd0; 1219: data <= 'd0; 1220: data <= 'd0; 1221: data <= 'd0; 1222: data <= 'd0; 1223: data <= 'd0; 1224: data <= 'd0; 1225: data <= 'd0; 1226: data <= 'd0; 1227: data <= 'd0; 1228: data <= 'd0; 1229: data <= 'd0; 1230: data <= 'd0; 1231: data <= 'd0; 1232: data <= 'd0; 1233: data <= 'd0; 1234: data <= 'd0; 1235: data <= 'd0; 1236: data <= 'd0; 1237: data <= 'd0; 1238: data <= 'd0; 1239: data <= 'd0; 1240: data <= 'd0; 1241: data <= 'd0; 1242: data <= 'd0; 1243: data <= 'd0; 1244: data <= 'd0; 1245: data <= 'd0; 1246: data <= 'd0; 1247: data <= 'd0; 1248: data <= 'd0; 1249: data <= 'd0; 1250: data <= 'd0; 1251: data <= 'd0; 1252: data <= 'd0; 1253: data <= 'd0; 1254: data <= 'd0; 1255: data <= 'd0; 1256: data <= 'd0; 1257: data <= 'd0; 1258: data <= 'd0; 1259: data <= 'd0; 1260: data <= 'd0; 1261: data <= 'd0; 1262: data <= 'd0; 1263: data <= 'd0; 1264: data <= 'd0; 1265: data <= 'd0; 1266: data <= 'd0; 1267: data <= 'd0; 1268: data <= 'd0; 1269: data <= 'd0; 1270: data <= 'd0; 1271: data <= 'd0; 1272: data <= 'd0; 1273: data <= 'd0; 1274: data <= 'd0; 1275: data <= 'd1; 1276: data <= 'd1; 1277: data <= 'd1; 1278: data <= 'd1; 1279: data <= 'd1; 1280: data <= 'd0; 1281: data <= 'd0; 1282: data <= 'd0; 1283: data <= 'd0; 1284: data <= 'd0; 1285: data <= 'd0; 1286: data <= 'd0; 1287: data <= 'd0; 1288: data <= 'd0; 1289: data <= 'd0; 1290: data <= 'd0; 1291: data <= 'd0; 1292: data <= 'd0; 1293: data <= 'd0; 1294: data <= 'd0; 1295: data <= 'd0; 1296: data <= 'd0; 1297: data <= 'd0; 1298: data <= 'd0; 1299: data <= 'd1; 1300: data <= 'd1; 1301: data <= 'd1; 1302: data <= 'd1; 1303: data <= 'd1; 1304: data <= 'd1; 1305: data <= 'd1; 1306: data <= 'd1; 1307: data <= 'd1; 1308: data <= 'd0; 1309: data <= 'd0; 1310: data <= 'd0; 1311: data <= 'd0; 1312: data <= 'd0; 1313: data <= 'd0; 1314: data <= 'd0; 1315: data <= 'd0; 1316: data <= 'd0; 1317: data <= 'd0; 1318: data <= 'd0; 1319: data <= 'd0; 1320: data <= 'd0; 1321: data <= 'd0; 1322: data <= 'd0; 1323: data <= 'd0; 1324: data <= 'd0; 1325: data <= 'd0; 1326: data <= 'd0; 1327: data <= 'd0; 1328: data <= 'd0; 1329: data <= 'd0; 1330: data <= 'd0; 1331: data <= 'd0; 1332: data <= 'd0; 1333: data <= 'd0; 1334: data <= 'd0; 1335: data <= 'd0; 1336: data <= 'd0; 1337: data <= 'd0; 1338: data <= 'd0; 1339: data <= 'd0; 1340: data <= 'd0; 1341: data <= 'd0; 1342: data <= 'd0; 1343: data <= 'd0; 1344: data <= 'd0; 1345: data <= 'd0; 1346: data <= 'd0; 1347: data <= 'd0; 1348: data <= 'd0; 1349: data <= 'd0; 1350: data <= 'd0; 1351: data <= 'd0; 1352: data <= 'd0; 1353: data <= 'd0; 1354: data <= 'd0; 1355: data <= 'd0; 1356: data <= 'd0; 1357: data <= 'd0; 1358: data <= 'd0; 1359: data <= 'd0; 1360: data <= 'd0; 1361: data <= 'd0; 1362: data <= 'd0; 1363: data <= 'd0; 1364: data <= 'd0; 1365: data <= 'd0; 1366: data <= 'd0; 1367: data <= 'd0; 1368: data <= 'd0; 1369: data <= 'd0; 1370: data <= 'd0; 1371: data <= 'd0; 1372: data <= 'd0; 1373: data <= 'd0; 1374: data <= 'd0; 1375: data <= 'd0; 1376: data <= 'd0; 1377: data <= 'd0; 1378: data <= 'd0; 1379: data <= 'd0; 1380: data <= 'd0; 1381: data <= 'd0; 1382: data <= 'd0; 1383: data <= 'd0; 1384: data <= 'd0; 1385: data <= 'd0; 1386: data <= 'd0; 1387: data <= 'd0; 1388: data <= 'd0; 1389: data <= 'd0; 1390: data <= 'd0; 1391: data <= 'd0; 1392: data <= 'd0; 1393: data <= 'd0; 1394: data <= 'd0; 1395: data <= 'd0; 1396: data <= 'd0; 1397: data <= 'd0; 1398: data <= 'd0; 1399: data <= 'd0; 1400: data <= 'd0; 1401: data <= 'd0; 1402: data <= 'd1; 1403: data <= 'd1; 1404: data <= 'd1; 1405: data <= 'd1; 1406: data <= 'd1; 1407: data <= 'd1; 1408: data <= 'd0; 1409: data <= 'd0; 1410: data <= 'd0; 1411: data <= 'd0; 1412: data <= 'd0; 1413: data <= 'd0; 1414: data <= 'd0; 1415: data <= 'd0; 1416: data <= 'd0; 1417: data <= 'd0; 1418: data <= 'd0; 1419: data <= 'd0; 1420: data <= 'd0; 1421: data <= 'd0; 1422: data <= 'd0; 1423: data <= 'd0; 1424: data <= 'd0; 1425: data <= 'd0; 1426: data <= 'd1; 1427: data <= 'd1; 1428: data <= 'd0; 1429: data <= 'd0; 1430: data <= 'd0; 1431: data <= 'd1; 1432: data <= 'd1; 1433: data <= 'd1; 1434: data <= 'd1; 1435: data <= 'd1; 1436: data <= 'd1; 1437: data <= 'd0; 1438: data <= 'd0; 1439: data <= 'd0; 1440: data <= 'd0; 1441: data <= 'd0; 1442: data <= 'd0; 1443: data <= 'd0; 1444: data <= 'd1; 1445: data <= 'd1; 1446: data <= 'd1; 1447: data <= 'd1; 1448: data <= 'd1; 1449: data <= 'd0; 1450: data <= 'd0; 1451: data <= 'd0; 1452: data <= 'd0; 1453: data <= 'd0; 1454: data <= 'd0; 1455: data <= 'd0; 1456: data <= 'd0; 1457: data <= 'd0; 1458: data <= 'd0; 1459: data <= 'd0; 1460: data <= 'd0; 1461: data <= 'd0; 1462: data <= 'd0; 1463: data <= 'd0; 1464: data <= 'd0; 1465: data <= 'd0; 1466: data <= 'd0; 1467: data <= 'd0; 1468: data <= 'd0; 1469: data <= 'd0; 1470: data <= 'd0; 1471: data <= 'd0; 1472: data <= 'd0; 1473: data <= 'd0; 1474: data <= 'd0; 1475: data <= 'd0; 1476: data <= 'd0; 1477: data <= 'd0; 1478: data <= 'd0; 1479: data <= 'd0; 1480: data <= 'd0; 1481: data <= 'd0; 1482: data <= 'd0; 1483: data <= 'd0; 1484: data <= 'd0; 1485: data <= 'd0; 1486: data <= 'd0; 1487: data <= 'd0; 1488: data <= 'd0; 1489: data <= 'd0; 1490: data <= 'd0; 1491: data <= 'd0; 1492: data <= 'd0; 1493: data <= 'd0; 1494: data <= 'd0; 1495: data <= 'd0; 1496: data <= 'd0; 1497: data <= 'd0; 1498: data <= 'd0; 1499: data <= 'd0; 1500: data <= 'd0; 1501: data <= 'd0; 1502: data <= 'd0; 1503: data <= 'd0; 1504: data <= 'd0; 1505: data <= 'd0; 1506: data <= 'd0; 1507: data <= 'd0; 1508: data <= 'd0; 1509: data <= 'd0; 1510: data <= 'd0; 1511: data <= 'd0; 1512: data <= 'd0; 1513: data <= 'd0; 1514: data <= 'd0; 1515: data <= 'd0; 1516: data <= 'd0; 1517: data <= 'd0; 1518: data <= 'd0; 1519: data <= 'd0; 1520: data <= 'd0; 1521: data <= 'd0; 1522: data <= 'd0; 1523: data <= 'd0; 1524: data <= 'd0; 1525: data <= 'd0; 1526: data <= 'd0; 1527: data <= 'd0; 1528: data <= 'd0; 1529: data <= 'd1; 1530: data <= 'd1; 1531: data <= 'd1; 1532: data <= 'd1; 1533: data <= 'd1; 1534: data <= 'd1; 1535: data <= 'd1; 1536: data <= 'd0; 1537: data <= 'd0; 1538: data <= 'd0; 1539: data <= 'd0; 1540: data <= 'd0; 1541: data <= 'd0; 1542: data <= 'd0; 1543: data <= 'd0; 1544: data <= 'd0; 1545: data <= 'd0; 1546: data <= 'd0; 1547: data <= 'd0; 1548: data <= 'd0; 1549: data <= 'd0; 1550: data <= 'd0; 1551: data <= 'd0; 1552: data <= 'd0; 1553: data <= 'd0; 1554: data <= 'd1; 1555: data <= 'd0; 1556: data <= 'd0; 1557: data <= 'd0; 1558: data <= 'd0; 1559: data <= 'd0; 1560: data <= 'd0; 1561: data <= 'd0; 1562: data <= 'd1; 1563: data <= 'd1; 1564: data <= 'd1; 1565: data <= 'd1; 1566: data <= 'd1; 1567: data <= 'd1; 1568: data <= 'd1; 1569: data <= 'd1; 1570: data <= 'd1; 1571: data <= 'd1; 1572: data <= 'd1; 1573: data <= 'd1; 1574: data <= 'd1; 1575: data <= 'd1; 1576: data <= 'd1; 1577: data <= 'd1; 1578: data <= 'd1; 1579: data <= 'd1; 1580: data <= 'd0; 1581: data <= 'd0; 1582: data <= 'd0; 1583: data <= 'd0; 1584: data <= 'd0; 1585: data <= 'd0; 1586: data <= 'd0; 1587: data <= 'd0; 1588: data <= 'd0; 1589: data <= 'd0; 1590: data <= 'd0; 1591: data <= 'd0; 1592: data <= 'd0; 1593: data <= 'd0; 1594: data <= 'd0; 1595: data <= 'd0; 1596: data <= 'd0; 1597: data <= 'd0; 1598: data <= 'd0; 1599: data <= 'd0; 1600: data <= 'd0; 1601: data <= 'd0; 1602: data <= 'd0; 1603: data <= 'd0; 1604: data <= 'd0; 1605: data <= 'd0; 1606: data <= 'd0; 1607: data <= 'd0; 1608: data <= 'd0; 1609: data <= 'd0; 1610: data <= 'd0; 1611: data <= 'd0; 1612: data <= 'd0; 1613: data <= 'd0; 1614: data <= 'd0; 1615: data <= 'd0; 1616: data <= 'd0; 1617: data <= 'd0; 1618: data <= 'd0; 1619: data <= 'd0; 1620: data <= 'd0; 1621: data <= 'd0; 1622: data <= 'd0; 1623: data <= 'd0; 1624: data <= 'd0; 1625: data <= 'd0; 1626: data <= 'd0; 1627: data <= 'd0; 1628: data <= 'd0; 1629: data <= 'd0; 1630: data <= 'd0; 1631: data <= 'd0; 1632: data <= 'd0; 1633: data <= 'd0; 1634: data <= 'd0; 1635: data <= 'd0; 1636: data <= 'd0; 1637: data <= 'd0; 1638: data <= 'd0; 1639: data <= 'd0; 1640: data <= 'd0; 1641: data <= 'd0; 1642: data <= 'd0; 1643: data <= 'd0; 1644: data <= 'd0; 1645: data <= 'd0; 1646: data <= 'd0; 1647: data <= 'd0; 1648: data <= 'd0; 1649: data <= 'd0; 1650: data <= 'd0; 1651: data <= 'd0; 1652: data <= 'd0; 1653: data <= 'd0; 1654: data <= 'd0; 1655: data <= 'd0; 1656: data <= 'd1; 1657: data <= 'd1; 1658: data <= 'd1; 1659: data <= 'd1; 1660: data <= 'd1; 1661: data <= 'd1; 1662: data <= 'd1; 1663: data <= 'd1; 1664: data <= 'd0; 1665: data <= 'd0; 1666: data <= 'd0; 1667: data <= 'd0; 1668: data <= 'd0; 1669: data <= 'd0; 1670: data <= 'd0; 1671: data <= 'd0; 1672: data <= 'd0; 1673: data <= 'd0; 1674: data <= 'd0; 1675: data <= 'd0; 1676: data <= 'd0; 1677: data <= 'd0; 1678: data <= 'd0; 1679: data <= 'd0; 1680: data <= 'd0; 1681: data <= 'd0; 1682: data <= 'd0; 1683: data <= 'd0; 1684: data <= 'd0; 1685: data <= 'd0; 1686: data <= 'd0; 1687: data <= 'd0; 1688: data <= 'd0; 1689: data <= 'd0; 1690: data <= 'd1; 1691: data <= 'd1; 1692: data <= 'd1; 1693: data <= 'd1; 1694: data <= 'd1; 1695: data <= 'd1; 1696: data <= 'd1; 1697: data <= 'd1; 1698: data <= 'd1; 1699: data <= 'd1; 1700: data <= 'd1; 1701: data <= 'd1; 1702: data <= 'd1; 1703: data <= 'd1; 1704: data <= 'd1; 1705: data <= 'd1; 1706: data <= 'd1; 1707: data <= 'd1; 1708: data <= 'd1; 1709: data <= 'd0; 1710: data <= 'd0; 1711: data <= 'd0; 1712: data <= 'd0; 1713: data <= 'd0; 1714: data <= 'd0; 1715: data <= 'd0; 1716: data <= 'd0; 1717: data <= 'd0; 1718: data <= 'd0; 1719: data <= 'd0; 1720: data <= 'd0; 1721: data <= 'd0; 1722: data <= 'd0; 1723: data <= 'd0; 1724: data <= 'd0; 1725: data <= 'd0; 1726: data <= 'd0; 1727: data <= 'd0; 1728: data <= 'd0; 1729: data <= 'd0; 1730: data <= 'd0; 1731: data <= 'd0; 1732: data <= 'd0; 1733: data <= 'd0; 1734: data <= 'd0; 1735: data <= 'd0; 1736: data <= 'd0; 1737: data <= 'd0; 1738: data <= 'd0; 1739: data <= 'd0; 1740: data <= 'd0; 1741: data <= 'd0; 1742: data <= 'd0; 1743: data <= 'd1; 1744: data <= 'd1; 1745: data <= 'd1; 1746: data <= 'd1; 1747: data <= 'd1; 1748: data <= 'd0; 1749: data <= 'd0; 1750: data <= 'd0; 1751: data <= 'd0; 1752: data <= 'd0; 1753: data <= 'd0; 1754: data <= 'd0; 1755: data <= 'd0; 1756: data <= 'd0; 1757: data <= 'd0; 1758: data <= 'd0; 1759: data <= 'd0; 1760: data <= 'd0; 1761: data <= 'd0; 1762: data <= 'd0; 1763: data <= 'd0; 1764: data <= 'd0; 1765: data <= 'd0; 1766: data <= 'd0; 1767: data <= 'd0; 1768: data <= 'd0; 1769: data <= 'd0; 1770: data <= 'd0; 1771: data <= 'd0; 1772: data <= 'd0; 1773: data <= 'd0; 1774: data <= 'd0; 1775: data <= 'd0; 1776: data <= 'd0; 1777: data <= 'd0; 1778: data <= 'd0; 1779: data <= 'd0; 1780: data <= 'd0; 1781: data <= 'd0; 1782: data <= 'd1; 1783: data <= 'd1; 1784: data <= 'd1; 1785: data <= 'd1; 1786: data <= 'd1; 1787: data <= 'd1; 1788: data <= 'd1; 1789: data <= 'd1; 1790: data <= 'd1; 1791: data <= 'd1; 1792: data <= 'd0; 1793: data <= 'd0; 1794: data <= 'd0; 1795: data <= 'd0; 1796: data <= 'd0; 1797: data <= 'd0; 1798: data <= 'd0; 1799: data <= 'd0; 1800: data <= 'd0; 1801: data <= 'd0; 1802: data <= 'd0; 1803: data <= 'd0; 1804: data <= 'd0; 1805: data <= 'd0; 1806: data <= 'd0; 1807: data <= 'd0; 1808: data <= 'd0; 1809: data <= 'd0; 1810: data <= 'd0; 1811: data <= 'd0; 1812: data <= 'd0; 1813: data <= 'd0; 1814: data <= 'd0; 1815: data <= 'd0; 1816: data <= 'd0; 1817: data <= 'd0; 1818: data <= 'd0; 1819: data <= 'd1; 1820: data <= 'd1; 1821: data <= 'd1; 1822: data <= 'd1; 1823: data <= 'd1; 1824: data <= 'd1; 1825: data <= 'd1; 1826: data <= 'd1; 1827: data <= 'd1; 1828: data <= 'd1; 1829: data <= 'd1; 1830: data <= 'd1; 1831: data <= 'd1; 1832: data <= 'd1; 1833: data <= 'd1; 1834: data <= 'd1; 1835: data <= 'd1; 1836: data <= 'd1; 1837: data <= 'd1; 1838: data <= 'd0; 1839: data <= 'd0; 1840: data <= 'd0; 1841: data <= 'd0; 1842: data <= 'd0; 1843: data <= 'd0; 1844: data <= 'd0; 1845: data <= 'd0; 1846: data <= 'd0; 1847: data <= 'd0; 1848: data <= 'd0; 1849: data <= 'd0; 1850: data <= 'd0; 1851: data <= 'd0; 1852: data <= 'd0; 1853: data <= 'd0; 1854: data <= 'd0; 1855: data <= 'd0; 1856: data <= 'd0; 1857: data <= 'd0; 1858: data <= 'd0; 1859: data <= 'd0; 1860: data <= 'd0; 1861: data <= 'd0; 1862: data <= 'd0; 1863: data <= 'd0; 1864: data <= 'd0; 1865: data <= 'd0; 1866: data <= 'd0; 1867: data <= 'd0; 1868: data <= 'd0; 1869: data <= 'd0; 1870: data <= 'd1; 1871: data <= 'd1; 1872: data <= 'd1; 1873: data <= 'd1; 1874: data <= 'd1; 1875: data <= 'd1; 1876: data <= 'd1; 1877: data <= 'd0; 1878: data <= 'd0; 1879: data <= 'd0; 1880: data <= 'd0; 1881: data <= 'd0; 1882: data <= 'd1; 1883: data <= 'd1; 1884: data <= 'd1; 1885: data <= 'd1; 1886: data <= 'd1; 1887: data <= 'd1; 1888: data <= 'd1; 1889: data <= 'd1; 1890: data <= 'd1; 1891: data <= 'd1; 1892: data <= 'd1; 1893: data <= 'd1; 1894: data <= 'd0; 1895: data <= 'd0; 1896: data <= 'd0; 1897: data <= 'd0; 1898: data <= 'd0; 1899: data <= 'd0; 1900: data <= 'd0; 1901: data <= 'd0; 1902: data <= 'd0; 1903: data <= 'd0; 1904: data <= 'd0; 1905: data <= 'd0; 1906: data <= 'd1; 1907: data <= 'd1; 1908: data <= 'd1; 1909: data <= 'd1; 1910: data <= 'd1; 1911: data <= 'd1; 1912: data <= 'd1; 1913: data <= 'd1; 1914: data <= 'd1; 1915: data <= 'd1; 1916: data <= 'd1; 1917: data <= 'd1; 1918: data <= 'd1; 1919: data <= 'd1; 1920: data <= 'd0; 1921: data <= 'd0; 1922: data <= 'd0; 1923: data <= 'd0; 1924: data <= 'd0; 1925: data <= 'd0; 1926: data <= 'd0; 1927: data <= 'd0; 1928: data <= 'd0; 1929: data <= 'd0; 1930: data <= 'd0; 1931: data <= 'd0; 1932: data <= 'd0; 1933: data <= 'd0; 1934: data <= 'd0; 1935: data <= 'd0; 1936: data <= 'd0; 1937: data <= 'd0; 1938: data <= 'd0; 1939: data <= 'd0; 1940: data <= 'd0; 1941: data <= 'd0; 1942: data <= 'd0; 1943: data <= 'd0; 1944: data <= 'd0; 1945: data <= 'd0; 1946: data <= 'd0; 1947: data <= 'd0; 1948: data <= 'd1; 1949: data <= 'd1; 1950: data <= 'd1; 1951: data <= 'd1; 1952: data <= 'd1; 1953: data <= 'd1; 1954: data <= 'd1; 1955: data <= 'd1; 1956: data <= 'd1; 1957: data <= 'd1; 1958: data <= 'd1; 1959: data <= 'd1; 1960: data <= 'd1; 1961: data <= 'd1; 1962: data <= 'd1; 1963: data <= 'd1; 1964: data <= 'd1; 1965: data <= 'd1; 1966: data <= 'd1; 1967: data <= 'd0; 1968: data <= 'd0; 1969: data <= 'd0; 1970: data <= 'd0; 1971: data <= 'd0; 1972: data <= 'd0; 1973: data <= 'd0; 1974: data <= 'd0; 1975: data <= 'd0; 1976: data <= 'd0; 1977: data <= 'd0; 1978: data <= 'd0; 1979: data <= 'd0; 1980: data <= 'd0; 1981: data <= 'd0; 1982: data <= 'd0; 1983: data <= 'd0; 1984: data <= 'd0; 1985: data <= 'd0; 1986: data <= 'd0; 1987: data <= 'd0; 1988: data <= 'd0; 1989: data <= 'd0; 1990: data <= 'd0; 1991: data <= 'd0; 1992: data <= 'd0; 1993: data <= 'd0; 1994: data <= 'd0; 1995: data <= 'd0; 1996: data <= 'd0; 1997: data <= 'd1; 1998: data <= 'd1; 1999: data <= 'd1; 2000: data <= 'd1; 2001: data <= 'd1; 2002: data <= 'd1; 2003: data <= 'd1; 2004: data <= 'd1; 2005: data <= 'd1; 2006: data <= 'd1; 2007: data <= 'd1; 2008: data <= 'd1; 2009: data <= 'd1; 2010: data <= 'd1; 2011: data <= 'd1; 2012: data <= 'd1; 2013: data <= 'd1; 2014: data <= 'd1; 2015: data <= 'd1; 2016: data <= 'd1; 2017: data <= 'd1; 2018: data <= 'd1; 2019: data <= 'd1; 2020: data <= 'd1; 2021: data <= 'd1; 2022: data <= 'd1; 2023: data <= 'd1; 2024: data <= 'd1; 2025: data <= 'd1; 2026: data <= 'd1; 2027: data <= 'd1; 2028: data <= 'd1; 2029: data <= 'd1; 2030: data <= 'd1; 2031: data <= 'd1; 2032: data <= 'd1; 2033: data <= 'd1; 2034: data <= 'd1; 2035: data <= 'd1; 2036: data <= 'd1; 2037: data <= 'd1; 2038: data <= 'd1; 2039: data <= 'd1; 2040: data <= 'd1; 2041: data <= 'd1; 2042: data <= 'd1; 2043: data <= 'd1; 2044: data <= 'd1; 2045: data <= 'd1; 2046: data <= 'd1; 2047: data <= 'd1; 2048: data <= 'd0; 2049: data <= 'd0; 2050: data <= 'd0; 2051: data <= 'd0; 2052: data <= 'd0; 2053: data <= 'd0; 2054: data <= 'd0; 2055: data <= 'd0; 2056: data <= 'd0; 2057: data <= 'd0; 2058: data <= 'd0; 2059: data <= 'd0; 2060: data <= 'd0; 2061: data <= 'd0; 2062: data <= 'd0; 2063: data <= 'd0; 2064: data <= 'd0; 2065: data <= 'd0; 2066: data <= 'd0; 2067: data <= 'd0; 2068: data <= 'd0; 2069: data <= 'd0; 2070: data <= 'd0; 2071: data <= 'd0; 2072: data <= 'd0; 2073: data <= 'd0; 2074: data <= 'd0; 2075: data <= 'd0; 2076: data <= 'd0; 2077: data <= 'd0; 2078: data <= 'd0; 2079: data <= 'd0; 2080: data <= 'd0; 2081: data <= 'd0; 2082: data <= 'd1; 2083: data <= 'd1; 2084: data <= 'd1; 2085: data <= 'd1; 2086: data <= 'd1; 2087: data <= 'd1; 2088: data <= 'd1; 2089: data <= 'd1; 2090: data <= 'd1; 2091: data <= 'd1; 2092: data <= 'd1; 2093: data <= 'd1; 2094: data <= 'd1; 2095: data <= 'd1; 2096: data <= 'd0; 2097: data <= 'd0; 2098: data <= 'd0; 2099: data <= 'd0; 2100: data <= 'd0; 2101: data <= 'd0; 2102: data <= 'd0; 2103: data <= 'd0; 2104: data <= 'd0; 2105: data <= 'd0; 2106: data <= 'd0; 2107: data <= 'd0; 2108: data <= 'd0; 2109: data <= 'd0; 2110: data <= 'd0; 2111: data <= 'd0; 2112: data <= 'd0; 2113: data <= 'd0; 2114: data <= 'd0; 2115: data <= 'd0; 2116: data <= 'd0; 2117: data <= 'd0; 2118: data <= 'd0; 2119: data <= 'd0; 2120: data <= 'd0; 2121: data <= 'd0; 2122: data <= 'd0; 2123: data <= 'd0; 2124: data <= 'd1; 2125: data <= 'd1; 2126: data <= 'd1; 2127: data <= 'd1; 2128: data <= 'd1; 2129: data <= 'd1; 2130: data <= 'd1; 2131: data <= 'd1; 2132: data <= 'd1; 2133: data <= 'd1; 2134: data <= 'd1; 2135: data <= 'd1; 2136: data <= 'd1; 2137: data <= 'd1; 2138: data <= 'd1; 2139: data <= 'd1; 2140: data <= 'd1; 2141: data <= 'd1; 2142: data <= 'd1; 2143: data <= 'd1; 2144: data <= 'd1; 2145: data <= 'd1; 2146: data <= 'd1; 2147: data <= 'd1; 2148: data <= 'd1; 2149: data <= 'd1; 2150: data <= 'd1; 2151: data <= 'd1; 2152: data <= 'd1; 2153: data <= 'd1; 2154: data <= 'd1; 2155: data <= 'd1; 2156: data <= 'd1; 2157: data <= 'd1; 2158: data <= 'd1; 2159: data <= 'd1; 2160: data <= 'd1; 2161: data <= 'd1; 2162: data <= 'd1; 2163: data <= 'd1; 2164: data <= 'd1; 2165: data <= 'd1; 2166: data <= 'd1; 2167: data <= 'd1; 2168: data <= 'd1; 2169: data <= 'd1; 2170: data <= 'd1; 2171: data <= 'd1; 2172: data <= 'd1; 2173: data <= 'd1; 2174: data <= 'd1; 2175: data <= 'd1; 2176: data <= 'd0; 2177: data <= 'd0; 2178: data <= 'd0; 2179: data <= 'd0; 2180: data <= 'd0; 2181: data <= 'd0; 2182: data <= 'd0; 2183: data <= 'd0; 2184: data <= 'd0; 2185: data <= 'd0; 2186: data <= 'd0; 2187: data <= 'd0; 2188: data <= 'd0; 2189: data <= 'd0; 2190: data <= 'd0; 2191: data <= 'd0; 2192: data <= 'd0; 2193: data <= 'd0; 2194: data <= 'd0; 2195: data <= 'd0; 2196: data <= 'd0; 2197: data <= 'd0; 2198: data <= 'd0; 2199: data <= 'd0; 2200: data <= 'd0; 2201: data <= 'd0; 2202: data <= 'd0; 2203: data <= 'd0; 2204: data <= 'd0; 2205: data <= 'd0; 2206: data <= 'd0; 2207: data <= 'd1; 2208: data <= 'd1; 2209: data <= 'd1; 2210: data <= 'd1; 2211: data <= 'd1; 2212: data <= 'd1; 2213: data <= 'd1; 2214: data <= 'd1; 2215: data <= 'd1; 2216: data <= 'd1; 2217: data <= 'd1; 2218: data <= 'd1; 2219: data <= 'd1; 2220: data <= 'd1; 2221: data <= 'd1; 2222: data <= 'd1; 2223: data <= 'd1; 2224: data <= 'd1; 2225: data <= 'd1; 2226: data <= 'd1; 2227: data <= 'd1; 2228: data <= 'd1; 2229: data <= 'd1; 2230: data <= 'd1; 2231: data <= 'd1; 2232: data <= 'd1; 2233: data <= 'd1; 2234: data <= 'd0; 2235: data <= 'd0; 2236: data <= 'd0; 2237: data <= 'd0; 2238: data <= 'd0; 2239: data <= 'd0; 2240: data <= 'd0; 2241: data <= 'd0; 2242: data <= 'd0; 2243: data <= 'd0; 2244: data <= 'd0; 2245: data <= 'd0; 2246: data <= 'd0; 2247: data <= 'd0; 2248: data <= 'd1; 2249: data <= 'd1; 2250: data <= 'd1; 2251: data <= 'd1; 2252: data <= 'd1; 2253: data <= 'd1; 2254: data <= 'd1; 2255: data <= 'd1; 2256: data <= 'd1; 2257: data <= 'd1; 2258: data <= 'd1; 2259: data <= 'd1; 2260: data <= 'd1; 2261: data <= 'd1; 2262: data <= 'd1; 2263: data <= 'd1; 2264: data <= 'd1; 2265: data <= 'd1; 2266: data <= 'd1; 2267: data <= 'd1; 2268: data <= 'd1; 2269: data <= 'd1; 2270: data <= 'd1; 2271: data <= 'd1; 2272: data <= 'd1; 2273: data <= 'd1; 2274: data <= 'd1; 2275: data <= 'd1; 2276: data <= 'd1; 2277: data <= 'd1; 2278: data <= 'd1; 2279: data <= 'd1; 2280: data <= 'd1; 2281: data <= 'd1; 2282: data <= 'd1; 2283: data <= 'd1; 2284: data <= 'd1; 2285: data <= 'd1; 2286: data <= 'd1; 2287: data <= 'd1; 2288: data <= 'd1; 2289: data <= 'd1; 2290: data <= 'd1; 2291: data <= 'd1; 2292: data <= 'd1; 2293: data <= 'd1; 2294: data <= 'd1; 2295: data <= 'd1; 2296: data <= 'd1; 2297: data <= 'd1; 2298: data <= 'd1; 2299: data <= 'd1; 2300: data <= 'd1; 2301: data <= 'd1; 2302: data <= 'd1; 2303: data <= 'd1; 2304: data <= 'd0; 2305: data <= 'd0; 2306: data <= 'd0; 2307: data <= 'd0; 2308: data <= 'd0; 2309: data <= 'd0; 2310: data <= 'd0; 2311: data <= 'd1; 2312: data <= 'd1; 2313: data <= 'd1; 2314: data <= 'd1; 2315: data <= 'd0; 2316: data <= 'd0; 2317: data <= 'd0; 2318: data <= 'd0; 2319: data <= 'd0; 2320: data <= 'd0; 2321: data <= 'd0; 2322: data <= 'd0; 2323: data <= 'd0; 2324: data <= 'd0; 2325: data <= 'd0; 2326: data <= 'd0; 2327: data <= 'd0; 2328: data <= 'd0; 2329: data <= 'd0; 2330: data <= 'd0; 2331: data <= 'd0; 2332: data <= 'd1; 2333: data <= 'd1; 2334: data <= 'd1; 2335: data <= 'd1; 2336: data <= 'd1; 2337: data <= 'd1; 2338: data <= 'd1; 2339: data <= 'd1; 2340: data <= 'd1; 2341: data <= 'd1; 2342: data <= 'd1; 2343: data <= 'd1; 2344: data <= 'd1; 2345: data <= 'd1; 2346: data <= 'd1; 2347: data <= 'd1; 2348: data <= 'd1; 2349: data <= 'd1; 2350: data <= 'd1; 2351: data <= 'd1; 2352: data <= 'd1; 2353: data <= 'd1; 2354: data <= 'd1; 2355: data <= 'd1; 2356: data <= 'd1; 2357: data <= 'd1; 2358: data <= 'd1; 2359: data <= 'd1; 2360: data <= 'd1; 2361: data <= 'd1; 2362: data <= 'd1; 2363: data <= 'd1; 2364: data <= 'd1; 2365: data <= 'd1; 2366: data <= 'd1; 2367: data <= 'd1; 2368: data <= 'd1; 2369: data <= 'd1; 2370: data <= 'd1; 2371: data <= 'd1; 2372: data <= 'd1; 2373: data <= 'd1; 2374: data <= 'd1; 2375: data <= 'd1; 2376: data <= 'd1; 2377: data <= 'd1; 2378: data <= 'd1; 2379: data <= 'd1; 2380: data <= 'd1; 2381: data <= 'd1; 2382: data <= 'd1; 2383: data <= 'd1; 2384: data <= 'd1; 2385: data <= 'd1; 2386: data <= 'd1; 2387: data <= 'd1; 2388: data <= 'd1; 2389: data <= 'd1; 2390: data <= 'd1; 2391: data <= 'd1; 2392: data <= 'd1; 2393: data <= 'd1; 2394: data <= 'd1; 2395: data <= 'd1; 2396: data <= 'd1; 2397: data <= 'd1; 2398: data <= 'd1; 2399: data <= 'd1; 2400: data <= 'd1; 2401: data <= 'd1; 2402: data <= 'd1; 2403: data <= 'd1; 2404: data <= 'd1; 2405: data <= 'd1; 2406: data <= 'd1; 2407: data <= 'd1; 2408: data <= 'd1; 2409: data <= 'd1; 2410: data <= 'd1; 2411: data <= 'd1; 2412: data <= 'd1; 2413: data <= 'd1; 2414: data <= 'd1; 2415: data <= 'd1; 2416: data <= 'd1; 2417: data <= 'd1; 2418: data <= 'd1; 2419: data <= 'd1; 2420: data <= 'd1; 2421: data <= 'd1; 2422: data <= 'd1; 2423: data <= 'd1; 2424: data <= 'd1; 2425: data <= 'd1; 2426: data <= 'd1; 2427: data <= 'd1; 2428: data <= 'd1; 2429: data <= 'd1; 2430: data <= 'd1; 2431: data <= 'd1; 2432: data <= 'd0; 2433: data <= 'd0; 2434: data <= 'd0; 2435: data <= 'd0; 2436: data <= 'd0; 2437: data <= 'd0; 2438: data <= 'd0; 2439: data <= 'd1; 2440: data <= 'd1; 2441: data <= 'd1; 2442: data <= 'd1; 2443: data <= 'd1; 2444: data <= 'd1; 2445: data <= 'd1; 2446: data <= 'd1; 2447: data <= 'd0; 2448: data <= 'd0; 2449: data <= 'd0; 2450: data <= 'd0; 2451: data <= 'd0; 2452: data <= 'd0; 2453: data <= 'd0; 2454: data <= 'd0; 2455: data <= 'd0; 2456: data <= 'd0; 2457: data <= 'd0; 2458: data <= 'd1; 2459: data <= 'd1; 2460: data <= 'd1; 2461: data <= 'd1; 2462: data <= 'd1; 2463: data <= 'd1; 2464: data <= 'd1; 2465: data <= 'd1; 2466: data <= 'd1; 2467: data <= 'd1; 2468: data <= 'd1; 2469: data <= 'd1; 2470: data <= 'd1; 2471: data <= 'd1; 2472: data <= 'd1; 2473: data <= 'd1; 2474: data <= 'd1; 2475: data <= 'd1; 2476: data <= 'd1; 2477: data <= 'd1; 2478: data <= 'd1; 2479: data <= 'd1; 2480: data <= 'd1; 2481: data <= 'd1; 2482: data <= 'd1; 2483: data <= 'd1; 2484: data <= 'd1; 2485: data <= 'd1; 2486: data <= 'd1; 2487: data <= 'd1; 2488: data <= 'd1; 2489: data <= 'd1; 2490: data <= 'd1; 2491: data <= 'd1; 2492: data <= 'd1; 2493: data <= 'd1; 2494: data <= 'd1; 2495: data <= 'd1; 2496: data <= 'd1; 2497: data <= 'd1; 2498: data <= 'd1; 2499: data <= 'd1; 2500: data <= 'd1; 2501: data <= 'd1; 2502: data <= 'd1; 2503: data <= 'd1; 2504: data <= 'd1; 2505: data <= 'd1; 2506: data <= 'd1; 2507: data <= 'd1; 2508: data <= 'd1; 2509: data <= 'd1; 2510: data <= 'd1; 2511: data <= 'd1; 2512: data <= 'd1; 2513: data <= 'd1; 2514: data <= 'd1; 2515: data <= 'd1; 2516: data <= 'd1; 2517: data <= 'd1; 2518: data <= 'd1; 2519: data <= 'd1; 2520: data <= 'd1; 2521: data <= 'd1; 2522: data <= 'd1; 2523: data <= 'd1; 2524: data <= 'd1; 2525: data <= 'd1; 2526: data <= 'd1; 2527: data <= 'd1; 2528: data <= 'd1; 2529: data <= 'd1; 2530: data <= 'd1; 2531: data <= 'd1; 2532: data <= 'd1; 2533: data <= 'd1; 2534: data <= 'd1; 2535: data <= 'd1; 2536: data <= 'd1; 2537: data <= 'd1; 2538: data <= 'd1; 2539: data <= 'd1; 2540: data <= 'd1; 2541: data <= 'd1; 2542: data <= 'd1; 2543: data <= 'd1; 2544: data <= 'd1; 2545: data <= 'd1; 2546: data <= 'd1; 2547: data <= 'd1; 2548: data <= 'd1; 2549: data <= 'd1; 2550: data <= 'd1; 2551: data <= 'd1; 2552: data <= 'd1; 2553: data <= 'd1; 2554: data <= 'd1; 2555: data <= 'd1; 2556: data <= 'd1; 2557: data <= 'd1; 2558: data <= 'd1; 2559: data <= 'd1; 2560: data <= 'd0; 2561: data <= 'd0; 2562: data <= 'd0; 2563: data <= 'd0; 2564: data <= 'd0; 2565: data <= 'd1; 2566: data <= 'd1; 2567: data <= 'd1; 2568: data <= 'd1; 2569: data <= 'd1; 2570: data <= 'd1; 2571: data <= 'd1; 2572: data <= 'd1; 2573: data <= 'd1; 2574: data <= 'd1; 2575: data <= 'd1; 2576: data <= 'd0; 2577: data <= 'd0; 2578: data <= 'd0; 2579: data <= 'd0; 2580: data <= 'd0; 2581: data <= 'd0; 2582: data <= 'd0; 2583: data <= 'd0; 2584: data <= 'd0; 2585: data <= 'd1; 2586: data <= 'd1; 2587: data <= 'd1; 2588: data <= 'd1; 2589: data <= 'd1; 2590: data <= 'd1; 2591: data <= 'd1; 2592: data <= 'd1; 2593: data <= 'd1; 2594: data <= 'd1; 2595: data <= 'd1; 2596: data <= 'd1; 2597: data <= 'd1; 2598: data <= 'd1; 2599: data <= 'd1; 2600: data <= 'd1; 2601: data <= 'd1; 2602: data <= 'd1; 2603: data <= 'd1; 2604: data <= 'd1; 2605: data <= 'd1; 2606: data <= 'd1; 2607: data <= 'd1; 2608: data <= 'd1; 2609: data <= 'd1; 2610: data <= 'd1; 2611: data <= 'd1; 2612: data <= 'd1; 2613: data <= 'd1; 2614: data <= 'd1; 2615: data <= 'd1; 2616: data <= 'd1; 2617: data <= 'd1; 2618: data <= 'd1; 2619: data <= 'd1; 2620: data <= 'd1; 2621: data <= 'd1; 2622: data <= 'd1; 2623: data <= 'd1; 2624: data <= 'd1; 2625: data <= 'd1; 2626: data <= 'd1; 2627: data <= 'd1; 2628: data <= 'd1; 2629: data <= 'd1; 2630: data <= 'd1; 2631: data <= 'd1; 2632: data <= 'd1; 2633: data <= 'd1; 2634: data <= 'd1; 2635: data <= 'd1; 2636: data <= 'd1; 2637: data <= 'd1; 2638: data <= 'd1; 2639: data <= 'd1; 2640: data <= 'd1; 2641: data <= 'd1; 2642: data <= 'd1; 2643: data <= 'd1; 2644: data <= 'd1; 2645: data <= 'd1; 2646: data <= 'd1; 2647: data <= 'd1; 2648: data <= 'd1; 2649: data <= 'd1; 2650: data <= 'd1; 2651: data <= 'd1; 2652: data <= 'd1; 2653: data <= 'd1; 2654: data <= 'd1; 2655: data <= 'd1; 2656: data <= 'd1; 2657: data <= 'd1; 2658: data <= 'd1; 2659: data <= 'd1; 2660: data <= 'd1; 2661: data <= 'd1; 2662: data <= 'd1; 2663: data <= 'd1; 2664: data <= 'd1; 2665: data <= 'd1; 2666: data <= 'd1; 2667: data <= 'd1; 2668: data <= 'd1; 2669: data <= 'd1; 2670: data <= 'd1; 2671: data <= 'd1; 2672: data <= 'd1; 2673: data <= 'd1; 2674: data <= 'd1; 2675: data <= 'd1; 2676: data <= 'd1; 2677: data <= 'd1; 2678: data <= 'd1; 2679: data <= 'd1; 2680: data <= 'd1; 2681: data <= 'd1; 2682: data <= 'd1; 2683: data <= 'd1; 2684: data <= 'd1; 2685: data <= 'd1; 2686: data <= 'd1; 2687: data <= 'd1; 2688: data <= 'd0; 2689: data <= 'd0; 2690: data <= 'd0; 2691: data <= 'd0; 2692: data <= 'd1; 2693: data <= 'd1; 2694: data <= 'd1; 2695: data <= 'd1; 2696: data <= 'd1; 2697: data <= 'd1; 2698: data <= 'd1; 2699: data <= 'd1; 2700: data <= 'd1; 2701: data <= 'd1; 2702: data <= 'd1; 2703: data <= 'd1; 2704: data <= 'd1; 2705: data <= 'd0; 2706: data <= 'd0; 2707: data <= 'd0; 2708: data <= 'd0; 2709: data <= 'd0; 2710: data <= 'd0; 2711: data <= 'd0; 2712: data <= 'd0; 2713: data <= 'd1; 2714: data <= 'd1; 2715: data <= 'd1; 2716: data <= 'd1; 2717: data <= 'd1; 2718: data <= 'd1; 2719: data <= 'd1; 2720: data <= 'd1; 2721: data <= 'd1; 2722: data <= 'd1; 2723: data <= 'd1; 2724: data <= 'd1; 2725: data <= 'd1; 2726: data <= 'd1; 2727: data <= 'd1; 2728: data <= 'd1; 2729: data <= 'd1; 2730: data <= 'd1; 2731: data <= 'd1; 2732: data <= 'd1; 2733: data <= 'd1; 2734: data <= 'd1; 2735: data <= 'd1; 2736: data <= 'd1; 2737: data <= 'd1; 2738: data <= 'd1; 2739: data <= 'd1; 2740: data <= 'd1; 2741: data <= 'd1; 2742: data <= 'd1; 2743: data <= 'd1; 2744: data <= 'd1; 2745: data <= 'd1; 2746: data <= 'd1; 2747: data <= 'd1; 2748: data <= 'd1; 2749: data <= 'd1; 2750: data <= 'd1; 2751: data <= 'd1; 2752: data <= 'd1; 2753: data <= 'd1; 2754: data <= 'd1; 2755: data <= 'd1; 2756: data <= 'd1; 2757: data <= 'd1; 2758: data <= 'd1; 2759: data <= 'd1; 2760: data <= 'd1; 2761: data <= 'd1; 2762: data <= 'd1; 2763: data <= 'd1; 2764: data <= 'd1; 2765: data <= 'd1; 2766: data <= 'd1; 2767: data <= 'd1; 2768: data <= 'd1; 2769: data <= 'd1; 2770: data <= 'd1; 2771: data <= 'd1; 2772: data <= 'd1; 2773: data <= 'd1; 2774: data <= 'd1; 2775: data <= 'd1; 2776: data <= 'd1; 2777: data <= 'd1; 2778: data <= 'd1; 2779: data <= 'd1; 2780: data <= 'd1; 2781: data <= 'd1; 2782: data <= 'd1; 2783: data <= 'd1; 2784: data <= 'd1; 2785: data <= 'd1; 2786: data <= 'd1; 2787: data <= 'd1; 2788: data <= 'd1; 2789: data <= 'd1; 2790: data <= 'd1; 2791: data <= 'd1; 2792: data <= 'd1; 2793: data <= 'd1; 2794: data <= 'd1; 2795: data <= 'd1; 2796: data <= 'd1; 2797: data <= 'd1; 2798: data <= 'd1; 2799: data <= 'd1; 2800: data <= 'd1; 2801: data <= 'd1; 2802: data <= 'd1; 2803: data <= 'd1; 2804: data <= 'd1; 2805: data <= 'd1; 2806: data <= 'd1; 2807: data <= 'd1; 2808: data <= 'd1; 2809: data <= 'd1; 2810: data <= 'd1; 2811: data <= 'd1; 2812: data <= 'd1; 2813: data <= 'd1; 2814: data <= 'd1; 2815: data <= 'd1; 2816: data <= 'd0; 2817: data <= 'd0; 2818: data <= 'd0; 2819: data <= 'd0; 2820: data <= 'd1; 2821: data <= 'd1; 2822: data <= 'd1; 2823: data <= 'd1; 2824: data <= 'd1; 2825: data <= 'd1; 2826: data <= 'd1; 2827: data <= 'd1; 2828: data <= 'd1; 2829: data <= 'd1; 2830: data <= 'd1; 2831: data <= 'd1; 2832: data <= 'd1; 2833: data <= 'd1; 2834: data <= 'd0; 2835: data <= 'd0; 2836: data <= 'd0; 2837: data <= 'd0; 2838: data <= 'd0; 2839: data <= 'd0; 2840: data <= 'd1; 2841: data <= 'd1; 2842: data <= 'd1; 2843: data <= 'd1; 2844: data <= 'd1; 2845: data <= 'd1; 2846: data <= 'd1; 2847: data <= 'd1; 2848: data <= 'd1; 2849: data <= 'd1; 2850: data <= 'd1; 2851: data <= 'd1; 2852: data <= 'd1; 2853: data <= 'd1; 2854: data <= 'd1; 2855: data <= 'd1; 2856: data <= 'd1; 2857: data <= 'd1; 2858: data <= 'd1; 2859: data <= 'd1; 2860: data <= 'd1; 2861: data <= 'd1; 2862: data <= 'd1; 2863: data <= 'd1; 2864: data <= 'd1; 2865: data <= 'd1; 2866: data <= 'd1; 2867: data <= 'd1; 2868: data <= 'd1; 2869: data <= 'd1; 2870: data <= 'd1; 2871: data <= 'd1; 2872: data <= 'd1; 2873: data <= 'd1; 2874: data <= 'd1; 2875: data <= 'd1; 2876: data <= 'd1; 2877: data <= 'd1; 2878: data <= 'd1; 2879: data <= 'd1; 2880: data <= 'd1; 2881: data <= 'd1; 2882: data <= 'd1; 2883: data <= 'd1; 2884: data <= 'd1; 2885: data <= 'd1; 2886: data <= 'd1; 2887: data <= 'd1; 2888: data <= 'd1; 2889: data <= 'd1; 2890: data <= 'd1; 2891: data <= 'd1; 2892: data <= 'd1; 2893: data <= 'd1; 2894: data <= 'd1; 2895: data <= 'd1; 2896: data <= 'd1; 2897: data <= 'd1; 2898: data <= 'd1; 2899: data <= 'd1; 2900: data <= 'd1; 2901: data <= 'd1; 2902: data <= 'd1; 2903: data <= 'd1; 2904: data <= 'd1; 2905: data <= 'd1; 2906: data <= 'd1; 2907: data <= 'd1; 2908: data <= 'd1; 2909: data <= 'd1; 2910: data <= 'd1; 2911: data <= 'd1; 2912: data <= 'd1; 2913: data <= 'd1; 2914: data <= 'd1; 2915: data <= 'd1; 2916: data <= 'd1; 2917: data <= 'd1; 2918: data <= 'd1; 2919: data <= 'd1; 2920: data <= 'd1; 2921: data <= 'd1; 2922: data <= 'd1; 2923: data <= 'd1; 2924: data <= 'd1; 2925: data <= 'd1; 2926: data <= 'd1; 2927: data <= 'd1; 2928: data <= 'd1; 2929: data <= 'd1; 2930: data <= 'd1; 2931: data <= 'd1; 2932: data <= 'd1; 2933: data <= 'd1; 2934: data <= 'd1; 2935: data <= 'd1; 2936: data <= 'd1; 2937: data <= 'd1; 2938: data <= 'd1; 2939: data <= 'd1; 2940: data <= 'd1; 2941: data <= 'd1; 2942: data <= 'd1; 2943: data <= 'd1; 2944: data <= 'd0; 2945: data <= 'd0; 2946: data <= 'd0; 2947: data <= 'd1; 2948: data <= 'd1; 2949: data <= 'd1; 2950: data <= 'd1; 2951: data <= 'd1; 2952: data <= 'd1; 2953: data <= 'd1; 2954: data <= 'd1; 2955: data <= 'd1; 2956: data <= 'd1; 2957: data <= 'd1; 2958: data <= 'd1; 2959: data <= 'd1; 2960: data <= 'd1; 2961: data <= 'd1; 2962: data <= 'd1; 2963: data <= 'd1; 2964: data <= 'd1; 2965: data <= 'd1; 2966: data <= 'd1; 2967: data <= 'd1; 2968: data <= 'd1; 2969: data <= 'd1; 2970: data <= 'd1; 2971: data <= 'd1; 2972: data <= 'd1; 2973: data <= 'd1; 2974: data <= 'd1; 2975: data <= 'd1; 2976: data <= 'd1; 2977: data <= 'd1; 2978: data <= 'd1; 2979: data <= 'd1; 2980: data <= 'd1; 2981: data <= 'd1; 2982: data <= 'd1; 2983: data <= 'd1; 2984: data <= 'd1; 2985: data <= 'd1; 2986: data <= 'd1; 2987: data <= 'd1; 2988: data <= 'd1; 2989: data <= 'd1; 2990: data <= 'd1; 2991: data <= 'd1; 2992: data <= 'd1; 2993: data <= 'd1; 2994: data <= 'd1; 2995: data <= 'd1; 2996: data <= 'd1; 2997: data <= 'd1; 2998: data <= 'd1; 2999: data <= 'd1; 3000: data <= 'd1; 3001: data <= 'd1; 3002: data <= 'd1; 3003: data <= 'd1; 3004: data <= 'd1; 3005: data <= 'd1; 3006: data <= 'd1; 3007: data <= 'd1; 3008: data <= 'd1; 3009: data <= 'd1; 3010: data <= 'd1; 3011: data <= 'd1; 3012: data <= 'd1; 3013: data <= 'd1; 3014: data <= 'd1; 3015: data <= 'd1; 3016: data <= 'd1; 3017: data <= 'd1; 3018: data <= 'd1; 3019: data <= 'd1; 3020: data <= 'd1; 3021: data <= 'd1; 3022: data <= 'd1; 3023: data <= 'd1; 3024: data <= 'd1; 3025: data <= 'd1; 3026: data <= 'd1; 3027: data <= 'd1; 3028: data <= 'd1; 3029: data <= 'd1; 3030: data <= 'd1; 3031: data <= 'd1; 3032: data <= 'd1; 3033: data <= 'd1; 3034: data <= 'd1; 3035: data <= 'd1; 3036: data <= 'd1; 3037: data <= 'd1; 3038: data <= 'd1; 3039: data <= 'd1; 3040: data <= 'd1; 3041: data <= 'd1; 3042: data <= 'd1; 3043: data <= 'd1; 3044: data <= 'd1; 3045: data <= 'd1; 3046: data <= 'd1; 3047: data <= 'd1; 3048: data <= 'd1; 3049: data <= 'd1; 3050: data <= 'd1; 3051: data <= 'd1; 3052: data <= 'd1; 3053: data <= 'd1; 3054: data <= 'd1; 3055: data <= 'd1; 3056: data <= 'd1; 3057: data <= 'd1; 3058: data <= 'd1; 3059: data <= 'd1; 3060: data <= 'd1; 3061: data <= 'd1; 3062: data <= 'd1; 3063: data <= 'd1; 3064: data <= 'd1; 3065: data <= 'd1; 3066: data <= 'd1; 3067: data <= 'd1; 3068: data <= 'd1; 3069: data <= 'd1; 3070: data <= 'd1; 3071: data <= 'd1; 3072: data <= 'd0; 3073: data <= 'd0; 3074: data <= 'd0; 3075: data <= 'd1; 3076: data <= 'd1; 3077: data <= 'd1; 3078: data <= 'd1; 3079: data <= 'd1; 3080: data <= 'd1; 3081: data <= 'd1; 3082: data <= 'd1; 3083: data <= 'd1; 3084: data <= 'd1; 3085: data <= 'd1; 3086: data <= 'd1; 3087: data <= 'd1; 3088: data <= 'd1; 3089: data <= 'd1; 3090: data <= 'd1; 3091: data <= 'd1; 3092: data <= 'd1; 3093: data <= 'd1; 3094: data <= 'd1; 3095: data <= 'd1; 3096: data <= 'd1; 3097: data <= 'd1; 3098: data <= 'd1; 3099: data <= 'd1; 3100: data <= 'd1; 3101: data <= 'd1; 3102: data <= 'd1; 3103: data <= 'd1; 3104: data <= 'd1; 3105: data <= 'd1; 3106: data <= 'd1; 3107: data <= 'd1; 3108: data <= 'd1; 3109: data <= 'd1; 3110: data <= 'd1; 3111: data <= 'd1; 3112: data <= 'd1; 3113: data <= 'd1; 3114: data <= 'd1; 3115: data <= 'd1; 3116: data <= 'd1; 3117: data <= 'd1; 3118: data <= 'd1; 3119: data <= 'd1; 3120: data <= 'd1; 3121: data <= 'd1; 3122: data <= 'd1; 3123: data <= 'd1; 3124: data <= 'd1; 3125: data <= 'd1; 3126: data <= 'd1; 3127: data <= 'd1; 3128: data <= 'd1; 3129: data <= 'd1; 3130: data <= 'd1; 3131: data <= 'd1; 3132: data <= 'd1; 3133: data <= 'd1; 3134: data <= 'd1; 3135: data <= 'd1; 3136: data <= 'd1; 3137: data <= 'd1; 3138: data <= 'd1; 3139: data <= 'd1; 3140: data <= 'd1; 3141: data <= 'd1; 3142: data <= 'd1; 3143: data <= 'd1; 3144: data <= 'd1; 3145: data <= 'd1; 3146: data <= 'd1; 3147: data <= 'd1; 3148: data <= 'd1; 3149: data <= 'd1; 3150: data <= 'd1; 3151: data <= 'd1; 3152: data <= 'd1; 3153: data <= 'd1; 3154: data <= 'd1; 3155: data <= 'd1; 3156: data <= 'd1; 3157: data <= 'd1; 3158: data <= 'd1; 3159: data <= 'd1; 3160: data <= 'd1; 3161: data <= 'd1; 3162: data <= 'd1; 3163: data <= 'd1; 3164: data <= 'd1; 3165: data <= 'd1; 3166: data <= 'd1; 3167: data <= 'd1; 3168: data <= 'd1; 3169: data <= 'd1; 3170: data <= 'd1; 3171: data <= 'd1; 3172: data <= 'd1; 3173: data <= 'd1; 3174: data <= 'd1; 3175: data <= 'd1; 3176: data <= 'd1; 3177: data <= 'd1; 3178: data <= 'd1; 3179: data <= 'd1; 3180: data <= 'd1; 3181: data <= 'd1; 3182: data <= 'd1; 3183: data <= 'd1; 3184: data <= 'd1; 3185: data <= 'd1; 3186: data <= 'd1; 3187: data <= 'd1; 3188: data <= 'd1; 3189: data <= 'd1; 3190: data <= 'd1; 3191: data <= 'd1; 3192: data <= 'd1; 3193: data <= 'd1; 3194: data <= 'd1; 3195: data <= 'd1; 3196: data <= 'd1; 3197: data <= 'd1; 3198: data <= 'd1; 3199: data <= 'd1; 3200: data <= 'd0; 3201: data <= 'd0; 3202: data <= 'd1; 3203: data <= 'd1; 3204: data <= 'd1; 3205: data <= 'd1; 3206: data <= 'd1; 3207: data <= 'd1; 3208: data <= 'd1; 3209: data <= 'd1; 3210: data <= 'd1; 3211: data <= 'd1; 3212: data <= 'd1; 3213: data <= 'd1; 3214: data <= 'd1; 3215: data <= 'd1; 3216: data <= 'd1; 3217: data <= 'd1; 3218: data <= 'd1; 3219: data <= 'd1; 3220: data <= 'd1; 3221: data <= 'd1; 3222: data <= 'd1; 3223: data <= 'd1; 3224: data <= 'd1; 3225: data <= 'd1; 3226: data <= 'd1; 3227: data <= 'd1; 3228: data <= 'd1; 3229: data <= 'd1; 3230: data <= 'd1; 3231: data <= 'd1; 3232: data <= 'd1; 3233: data <= 'd1; 3234: data <= 'd1; 3235: data <= 'd1; 3236: data <= 'd1; 3237: data <= 'd1; 3238: data <= 'd1; 3239: data <= 'd1; 3240: data <= 'd1; 3241: data <= 'd1; 3242: data <= 'd1; 3243: data <= 'd1; 3244: data <= 'd1; 3245: data <= 'd1; 3246: data <= 'd1; 3247: data <= 'd1; 3248: data <= 'd1; 3249: data <= 'd1; 3250: data <= 'd1; 3251: data <= 'd1; 3252: data <= 'd1; 3253: data <= 'd1; 3254: data <= 'd1; 3255: data <= 'd1; 3256: data <= 'd1; 3257: data <= 'd1; 3258: data <= 'd1; 3259: data <= 'd1; 3260: data <= 'd1; 3261: data <= 'd1; 3262: data <= 'd1; 3263: data <= 'd1; 3264: data <= 'd1; 3265: data <= 'd1; 3266: data <= 'd1; 3267: data <= 'd1; 3268: data <= 'd1; 3269: data <= 'd1; 3270: data <= 'd1; 3271: data <= 'd1; 3272: data <= 'd1; 3273: data <= 'd1; 3274: data <= 'd1; 3275: data <= 'd1; 3276: data <= 'd1; 3277: data <= 'd1; 3278: data <= 'd1; 3279: data <= 'd1; 3280: data <= 'd1; 3281: data <= 'd1; 3282: data <= 'd1; 3283: data <= 'd1; 3284: data <= 'd1; 3285: data <= 'd1; 3286: data <= 'd1; 3287: data <= 'd1; 3288: data <= 'd1; 3289: data <= 'd1; 3290: data <= 'd1; 3291: data <= 'd1; 3292: data <= 'd1; 3293: data <= 'd1; 3294: data <= 'd1; 3295: data <= 'd1; 3296: data <= 'd1; 3297: data <= 'd1; 3298: data <= 'd1; 3299: data <= 'd1; 3300: data <= 'd1; 3301: data <= 'd1; 3302: data <= 'd1; 3303: data <= 'd1; 3304: data <= 'd1; 3305: data <= 'd1; 3306: data <= 'd1; 3307: data <= 'd1; 3308: data <= 'd1; 3309: data <= 'd1; 3310: data <= 'd1; 3311: data <= 'd1; 3312: data <= 'd1; 3313: data <= 'd1; 3314: data <= 'd1; 3315: data <= 'd1; 3316: data <= 'd1; 3317: data <= 'd1; 3318: data <= 'd1; 3319: data <= 'd1; 3320: data <= 'd1; 3321: data <= 'd1; 3322: data <= 'd1; 3323: data <= 'd1; 3324: data <= 'd1; 3325: data <= 'd1; 3326: data <= 'd1; 3327: data <= 'd1; 3328: data <= 'd0; 3329: data <= 'd0; 3330: data <= 'd1; 3331: data <= 'd1; 3332: data <= 'd1; 3333: data <= 'd1; 3334: data <= 'd1; 3335: data <= 'd1; 3336: data <= 'd1; 3337: data <= 'd1; 3338: data <= 'd1; 3339: data <= 'd1; 3340: data <= 'd1; 3341: data <= 'd1; 3342: data <= 'd1; 3343: data <= 'd1; 3344: data <= 'd1; 3345: data <= 'd1; 3346: data <= 'd1; 3347: data <= 'd1; 3348: data <= 'd1; 3349: data <= 'd1; 3350: data <= 'd1; 3351: data <= 'd1; 3352: data <= 'd1; 3353: data <= 'd1; 3354: data <= 'd1; 3355: data <= 'd1; 3356: data <= 'd1; 3357: data <= 'd1; 3358: data <= 'd1; 3359: data <= 'd1; 3360: data <= 'd1; 3361: data <= 'd1; 3362: data <= 'd1; 3363: data <= 'd1; 3364: data <= 'd1; 3365: data <= 'd1; 3366: data <= 'd1; 3367: data <= 'd1; 3368: data <= 'd1; 3369: data <= 'd1; 3370: data <= 'd1; 3371: data <= 'd1; 3372: data <= 'd1; 3373: data <= 'd1; 3374: data <= 'd1; 3375: data <= 'd1; 3376: data <= 'd1; 3377: data <= 'd1; 3378: data <= 'd1; 3379: data <= 'd1; 3380: data <= 'd1; 3381: data <= 'd1; 3382: data <= 'd1; 3383: data <= 'd1; 3384: data <= 'd1; 3385: data <= 'd1; 3386: data <= 'd1; 3387: data <= 'd1; 3388: data <= 'd1; 3389: data <= 'd1; 3390: data <= 'd1; 3391: data <= 'd1; 3392: data <= 'd1; 3393: data <= 'd1; 3394: data <= 'd1; 3395: data <= 'd1; 3396: data <= 'd1; 3397: data <= 'd1; 3398: data <= 'd1; 3399: data <= 'd1; 3400: data <= 'd1; 3401: data <= 'd1; 3402: data <= 'd1; 3403: data <= 'd1; 3404: data <= 'd1; 3405: data <= 'd1; 3406: data <= 'd1; 3407: data <= 'd1; 3408: data <= 'd1; 3409: data <= 'd1; 3410: data <= 'd1; 3411: data <= 'd1; 3412: data <= 'd1; 3413: data <= 'd1; 3414: data <= 'd1; 3415: data <= 'd1; 3416: data <= 'd1; 3417: data <= 'd1; 3418: data <= 'd1; 3419: data <= 'd1; 3420: data <= 'd1; 3421: data <= 'd1; 3422: data <= 'd1; 3423: data <= 'd1; 3424: data <= 'd1; 3425: data <= 'd1; 3426: data <= 'd1; 3427: data <= 'd1; 3428: data <= 'd1; 3429: data <= 'd1; 3430: data <= 'd1; 3431: data <= 'd1; 3432: data <= 'd1; 3433: data <= 'd1; 3434: data <= 'd1; 3435: data <= 'd1; 3436: data <= 'd1; 3437: data <= 'd1; 3438: data <= 'd1; 3439: data <= 'd1; 3440: data <= 'd1; 3441: data <= 'd1; 3442: data <= 'd1; 3443: data <= 'd1; 3444: data <= 'd1; 3445: data <= 'd1; 3446: data <= 'd1; 3447: data <= 'd1; 3448: data <= 'd1; 3449: data <= 'd1; 3450: data <= 'd1; 3451: data <= 'd1; 3452: data <= 'd1; 3453: data <= 'd1; 3454: data <= 'd1; 3455: data <= 'd1; 3456: data <= 'd0; 3457: data <= 'd1; 3458: data <= 'd1; 3459: data <= 'd1; 3460: data <= 'd1; 3461: data <= 'd1; 3462: data <= 'd1; 3463: data <= 'd1; 3464: data <= 'd1; 3465: data <= 'd1; 3466: data <= 'd1; 3467: data <= 'd1; 3468: data <= 'd1; 3469: data <= 'd1; 3470: data <= 'd1; 3471: data <= 'd1; 3472: data <= 'd1; 3473: data <= 'd1; 3474: data <= 'd1; 3475: data <= 'd1; 3476: data <= 'd1; 3477: data <= 'd1; 3478: data <= 'd1; 3479: data <= 'd1; 3480: data <= 'd1; 3481: data <= 'd1; 3482: data <= 'd1; 3483: data <= 'd1; 3484: data <= 'd1; 3485: data <= 'd1; 3486: data <= 'd1; 3487: data <= 'd1; 3488: data <= 'd1; 3489: data <= 'd1; 3490: data <= 'd1; 3491: data <= 'd1; 3492: data <= 'd1; 3493: data <= 'd1; 3494: data <= 'd0; 3495: data <= 'd0; 3496: data <= 'd0; 3497: data <= 'd0; 3498: data <= 'd0; 3499: data <= 'd0; 3500: data <= 'd0; 3501: data <= 'd0; 3502: data <= 'd1; 3503: data <= 'd1; 3504: data <= 'd1; 3505: data <= 'd1; 3506: data <= 'd1; 3507: data <= 'd1; 3508: data <= 'd1; 3509: data <= 'd1; 3510: data <= 'd1; 3511: data <= 'd1; 3512: data <= 'd1; 3513: data <= 'd1; 3514: data <= 'd1; 3515: data <= 'd1; 3516: data <= 'd1; 3517: data <= 'd1; 3518: data <= 'd1; 3519: data <= 'd1; 3520: data <= 'd1; 3521: data <= 'd1; 3522: data <= 'd1; 3523: data <= 'd1; 3524: data <= 'd1; 3525: data <= 'd1; 3526: data <= 'd1; 3527: data <= 'd1; 3528: data <= 'd1; 3529: data <= 'd1; 3530: data <= 'd1; 3531: data <= 'd1; 3532: data <= 'd1; 3533: data <= 'd1; 3534: data <= 'd1; 3535: data <= 'd1; 3536: data <= 'd1; 3537: data <= 'd1; 3538: data <= 'd1; 3539: data <= 'd1; 3540: data <= 'd1; 3541: data <= 'd1; 3542: data <= 'd1; 3543: data <= 'd1; 3544: data <= 'd1; 3545: data <= 'd1; 3546: data <= 'd1; 3547: data <= 'd1; 3548: data <= 'd1; 3549: data <= 'd1; 3550: data <= 'd1; 3551: data <= 'd1; 3552: data <= 'd1; 3553: data <= 'd1; 3554: data <= 'd1; 3555: data <= 'd1; 3556: data <= 'd1; 3557: data <= 'd1; 3558: data <= 'd1; 3559: data <= 'd1; 3560: data <= 'd1; 3561: data <= 'd1; 3562: data <= 'd1; 3563: data <= 'd1; 3564: data <= 'd1; 3565: data <= 'd1; 3566: data <= 'd1; 3567: data <= 'd1; 3568: data <= 'd1; 3569: data <= 'd1; 3570: data <= 'd1; 3571: data <= 'd1; 3572: data <= 'd1; 3573: data <= 'd1; 3574: data <= 'd1; 3575: data <= 'd1; 3576: data <= 'd1; 3577: data <= 'd1; 3578: data <= 'd1; 3579: data <= 'd1; 3580: data <= 'd1; 3581: data <= 'd1; 3582: data <= 'd1; 3583: data <= 'd1; 3584: data <= 'd0; 3585: data <= 'd1; 3586: data <= 'd1; 3587: data <= 'd1; 3588: data <= 'd1; 3589: data <= 'd1; 3590: data <= 'd1; 3591: data <= 'd1; 3592: data <= 'd1; 3593: data <= 'd1; 3594: data <= 'd1; 3595: data <= 'd1; 3596: data <= 'd1; 3597: data <= 'd1; 3598: data <= 'd1; 3599: data <= 'd1; 3600: data <= 'd1; 3601: data <= 'd1; 3602: data <= 'd1; 3603: data <= 'd1; 3604: data <= 'd1; 3605: data <= 'd1; 3606: data <= 'd1; 3607: data <= 'd1; 3608: data <= 'd1; 3609: data <= 'd1; 3610: data <= 'd1; 3611: data <= 'd1; 3612: data <= 'd1; 3613: data <= 'd1; 3614: data <= 'd1; 3615: data <= 'd1; 3616: data <= 'd1; 3617: data <= 'd1; 3618: data <= 'd1; 3619: data <= 'd1; 3620: data <= 'd0; 3621: data <= 'd0; 3622: data <= 'd0; 3623: data <= 'd0; 3624: data <= 'd0; 3625: data <= 'd0; 3626: data <= 'd0; 3627: data <= 'd0; 3628: data <= 'd0; 3629: data <= 'd0; 3630: data <= 'd0; 3631: data <= 'd0; 3632: data <= 'd1; 3633: data <= 'd1; 3634: data <= 'd1; 3635: data <= 'd1; 3636: data <= 'd1; 3637: data <= 'd1; 3638: data <= 'd1; 3639: data <= 'd1; 3640: data <= 'd1; 3641: data <= 'd1; 3642: data <= 'd1; 3643: data <= 'd1; 3644: data <= 'd1; 3645: data <= 'd1; 3646: data <= 'd1; 3647: data <= 'd1; 3648: data <= 'd1; 3649: data <= 'd1; 3650: data <= 'd1; 3651: data <= 'd1; 3652: data <= 'd1; 3653: data <= 'd1; 3654: data <= 'd1; 3655: data <= 'd1; 3656: data <= 'd1; 3657: data <= 'd1; 3658: data <= 'd1; 3659: data <= 'd1; 3660: data <= 'd1; 3661: data <= 'd1; 3662: data <= 'd1; 3663: data <= 'd1; 3664: data <= 'd1; 3665: data <= 'd1; 3666: data <= 'd1; 3667: data <= 'd1; 3668: data <= 'd1; 3669: data <= 'd1; 3670: data <= 'd1; 3671: data <= 'd1; 3672: data <= 'd1; 3673: data <= 'd1; 3674: data <= 'd1; 3675: data <= 'd1; 3676: data <= 'd1; 3677: data <= 'd1; 3678: data <= 'd1; 3679: data <= 'd1; 3680: data <= 'd1; 3681: data <= 'd1; 3682: data <= 'd1; 3683: data <= 'd1; 3684: data <= 'd1; 3685: data <= 'd1; 3686: data <= 'd1; 3687: data <= 'd1; 3688: data <= 'd1; 3689: data <= 'd1; 3690: data <= 'd1; 3691: data <= 'd1; 3692: data <= 'd1; 3693: data <= 'd1; 3694: data <= 'd1; 3695: data <= 'd1; 3696: data <= 'd1; 3697: data <= 'd1; 3698: data <= 'd1; 3699: data <= 'd1; 3700: data <= 'd1; 3701: data <= 'd1; 3702: data <= 'd1; 3703: data <= 'd1; 3704: data <= 'd1; 3705: data <= 'd1; 3706: data <= 'd1; 3707: data <= 'd1; 3708: data <= 'd1; 3709: data <= 'd1; 3710: data <= 'd1; 3711: data <= 'd1; 3712: data <= 'd0; 3713: data <= 'd1; 3714: data <= 'd1; 3715: data <= 'd1; 3716: data <= 'd1; 3717: data <= 'd1; 3718: data <= 'd0; 3719: data <= 'd0; 3720: data <= 'd0; 3721: data <= 'd0; 3722: data <= 'd0; 3723: data <= 'd0; 3724: data <= 'd0; 3725: data <= 'd1; 3726: data <= 'd1; 3727: data <= 'd1; 3728: data <= 'd1; 3729: data <= 'd1; 3730: data <= 'd1; 3731: data <= 'd1; 3732: data <= 'd1; 3733: data <= 'd1; 3734: data <= 'd1; 3735: data <= 'd1; 3736: data <= 'd1; 3737: data <= 'd1; 3738: data <= 'd1; 3739: data <= 'd1; 3740: data <= 'd1; 3741: data <= 'd1; 3742: data <= 'd1; 3743: data <= 'd1; 3744: data <= 'd1; 3745: data <= 'd1; 3746: data <= 'd1; 3747: data <= 'd0; 3748: data <= 'd0; 3749: data <= 'd0; 3750: data <= 'd0; 3751: data <= 'd0; 3752: data <= 'd0; 3753: data <= 'd0; 3754: data <= 'd0; 3755: data <= 'd0; 3756: data <= 'd0; 3757: data <= 'd0; 3758: data <= 'd0; 3759: data <= 'd0; 3760: data <= 'd0; 3761: data <= 'd0; 3762: data <= 'd1; 3763: data <= 'd1; 3764: data <= 'd1; 3765: data <= 'd1; 3766: data <= 'd1; 3767: data <= 'd1; 3768: data <= 'd1; 3769: data <= 'd1; 3770: data <= 'd1; 3771: data <= 'd1; 3772: data <= 'd1; 3773: data <= 'd1; 3774: data <= 'd1; 3775: data <= 'd1; 3776: data <= 'd1; 3777: data <= 'd1; 3778: data <= 'd1; 3779: data <= 'd1; 3780: data <= 'd1; 3781: data <= 'd1; 3782: data <= 'd1; 3783: data <= 'd1; 3784: data <= 'd1; 3785: data <= 'd1; 3786: data <= 'd1; 3787: data <= 'd1; 3788: data <= 'd1; 3789: data <= 'd1; 3790: data <= 'd1; 3791: data <= 'd1; 3792: data <= 'd1; 3793: data <= 'd1; 3794: data <= 'd1; 3795: data <= 'd1; 3796: data <= 'd1; 3797: data <= 'd1; 3798: data <= 'd1; 3799: data <= 'd1; 3800: data <= 'd1; 3801: data <= 'd1; 3802: data <= 'd1; 3803: data <= 'd1; 3804: data <= 'd1; 3805: data <= 'd1; 3806: data <= 'd1; 3807: data <= 'd1; 3808: data <= 'd1; 3809: data <= 'd1; 3810: data <= 'd1; 3811: data <= 'd1; 3812: data <= 'd1; 3813: data <= 'd1; 3814: data <= 'd1; 3815: data <= 'd1; 3816: data <= 'd1; 3817: data <= 'd1; 3818: data <= 'd1; 3819: data <= 'd1; 3820: data <= 'd1; 3821: data <= 'd1; 3822: data <= 'd1; 3823: data <= 'd1; 3824: data <= 'd1; 3825: data <= 'd1; 3826: data <= 'd1; 3827: data <= 'd1; 3828: data <= 'd1; 3829: data <= 'd1; 3830: data <= 'd1; 3831: data <= 'd1; 3832: data <= 'd1; 3833: data <= 'd1; 3834: data <= 'd1; 3835: data <= 'd1; 3836: data <= 'd1; 3837: data <= 'd1; 3838: data <= 'd1; 3839: data <= 'd1; 3840: data <= 'd1; 3841: data <= 'd1; 3842: data <= 'd1; 3843: data <= 'd1; 3844: data <= 'd0; 3845: data <= 'd0; 3846: data <= 'd0; 3847: data <= 'd0; 3848: data <= 'd0; 3849: data <= 'd0; 3850: data <= 'd0; 3851: data <= 'd0; 3852: data <= 'd0; 3853: data <= 'd1; 3854: data <= 'd1; 3855: data <= 'd1; 3856: data <= 'd1; 3857: data <= 'd1; 3858: data <= 'd1; 3859: data <= 'd1; 3860: data <= 'd1; 3861: data <= 'd1; 3862: data <= 'd1; 3863: data <= 'd1; 3864: data <= 'd1; 3865: data <= 'd1; 3866: data <= 'd1; 3867: data <= 'd1; 3868: data <= 'd1; 3869: data <= 'd1; 3870: data <= 'd1; 3871: data <= 'd1; 3872: data <= 'd1; 3873: data <= 'd0; 3874: data <= 'd0; 3875: data <= 'd0; 3876: data <= 'd0; 3877: data <= 'd0; 3878: data <= 'd0; 3879: data <= 'd0; 3880: data <= 'd0; 3881: data <= 'd0; 3882: data <= 'd0; 3883: data <= 'd0; 3884: data <= 'd0; 3885: data <= 'd0; 3886: data <= 'd0; 3887: data <= 'd0; 3888: data <= 'd0; 3889: data <= 'd0; 3890: data <= 'd0; 3891: data <= 'd0; 3892: data <= 'd1; 3893: data <= 'd1; 3894: data <= 'd1; 3895: data <= 'd1; 3896: data <= 'd1; 3897: data <= 'd1; 3898: data <= 'd1; 3899: data <= 'd1; 3900: data <= 'd1; 3901: data <= 'd1; 3902: data <= 'd1; 3903: data <= 'd1; 3904: data <= 'd1; 3905: data <= 'd1; 3906: data <= 'd1; 3907: data <= 'd1; 3908: data <= 'd1; 3909: data <= 'd1; 3910: data <= 'd1; 3911: data <= 'd1; 3912: data <= 'd1; 3913: data <= 'd1; 3914: data <= 'd1; 3915: data <= 'd1; 3916: data <= 'd1; 3917: data <= 'd1; 3918: data <= 'd1; 3919: data <= 'd1; 3920: data <= 'd1; 3921: data <= 'd1; 3922: data <= 'd1; 3923: data <= 'd1; 3924: data <= 'd1; 3925: data <= 'd1; 3926: data <= 'd1; 3927: data <= 'd1; 3928: data <= 'd1; 3929: data <= 'd1; 3930: data <= 'd0; 3931: data <= 'd0; 3932: data <= 'd0; 3933: data <= 'd0; 3934: data <= 'd0; 3935: data <= 'd0; 3936: data <= 'd0; 3937: data <= 'd0; 3938: data <= 'd0; 3939: data <= 'd0; 3940: data <= 'd0; 3941: data <= 'd0; 3942: data <= 'd0; 3943: data <= 'd0; 3944: data <= 'd1; 3945: data <= 'd1; 3946: data <= 'd1; 3947: data <= 'd1; 3948: data <= 'd1; 3949: data <= 'd1; 3950: data <= 'd1; 3951: data <= 'd1; 3952: data <= 'd1; 3953: data <= 'd1; 3954: data <= 'd1; 3955: data <= 'd1; 3956: data <= 'd1; 3957: data <= 'd1; 3958: data <= 'd1; 3959: data <= 'd1; 3960: data <= 'd1; 3961: data <= 'd1; 3962: data <= 'd1; 3963: data <= 'd1; 3964: data <= 'd1; 3965: data <= 'd1; 3966: data <= 'd1; 3967: data <= 'd1; 3968: data <= 'd1; 3969: data <= 'd1; 3970: data <= 'd1; 3971: data <= 'd0; 3972: data <= 'd0; 3973: data <= 'd0; 3974: data <= 'd0; 3975: data <= 'd0; 3976: data <= 'd0; 3977: data <= 'd0; 3978: data <= 'd0; 3979: data <= 'd0; 3980: data <= 'd0; 3981: data <= 'd1; 3982: data <= 'd1; 3983: data <= 'd1; 3984: data <= 'd1; 3985: data <= 'd1; 3986: data <= 'd1; 3987: data <= 'd1; 3988: data <= 'd1; 3989: data <= 'd1; 3990: data <= 'd1; 3991: data <= 'd1; 3992: data <= 'd1; 3993: data <= 'd1; 3994: data <= 'd1; 3995: data <= 'd1; 3996: data <= 'd1; 3997: data <= 'd1; 3998: data <= 'd1; 3999: data <= 'd0; 4000: data <= 'd0; 4001: data <= 'd0; 4002: data <= 'd0; 4003: data <= 'd0; 4004: data <= 'd0; 4005: data <= 'd0; 4006: data <= 'd0; 4007: data <= 'd0; 4008: data <= 'd0; 4009: data <= 'd0; 4010: data <= 'd0; 4011: data <= 'd0; 4012: data <= 'd0; 4013: data <= 'd0; 4014: data <= 'd0; 4015: data <= 'd0; 4016: data <= 'd0; 4017: data <= 'd0; 4018: data <= 'd0; 4019: data <= 'd0; 4020: data <= 'd0; 4021: data <= 'd0; 4022: data <= 'd0; 4023: data <= 'd0; 4024: data <= 'd0; 4025: data <= 'd1; 4026: data <= 'd1; 4027: data <= 'd1; 4028: data <= 'd1; 4029: data <= 'd1; 4030: data <= 'd1; 4031: data <= 'd1; 4032: data <= 'd1; 4033: data <= 'd1; 4034: data <= 'd1; 4035: data <= 'd1; 4036: data <= 'd1; 4037: data <= 'd1; 4038: data <= 'd1; 4039: data <= 'd1; 4040: data <= 'd1; 4041: data <= 'd1; 4042: data <= 'd1; 4043: data <= 'd1; 4044: data <= 'd1; 4045: data <= 'd1; 4046: data <= 'd1; 4047: data <= 'd1; 4048: data <= 'd1; 4049: data <= 'd1; 4050: data <= 'd1; 4051: data <= 'd0; 4052: data <= 'd0; 4053: data <= 'd0; 4054: data <= 'd0; 4055: data <= 'd0; 4056: data <= 'd0; 4057: data <= 'd0; 4058: data <= 'd0; 4059: data <= 'd0; 4060: data <= 'd0; 4061: data <= 'd0; 4062: data <= 'd0; 4063: data <= 'd0; 4064: data <= 'd0; 4065: data <= 'd0; 4066: data <= 'd0; 4067: data <= 'd0; 4068: data <= 'd0; 4069: data <= 'd0; 4070: data <= 'd0; 4071: data <= 'd0; 4072: data <= 'd0; 4073: data <= 'd1; 4074: data <= 'd1; 4075: data <= 'd1; 4076: data <= 'd1; 4077: data <= 'd1; 4078: data <= 'd1; 4079: data <= 'd1; 4080: data <= 'd1; 4081: data <= 'd1; 4082: data <= 'd1; 4083: data <= 'd1; 4084: data <= 'd1; 4085: data <= 'd1; 4086: data <= 'd1; 4087: data <= 'd1; 4088: data <= 'd1; 4089: data <= 'd1; 4090: data <= 'd1; 4091: data <= 'd1; 4092: data <= 'd1; 4093: data <= 'd1; 4094: data <= 'd1; 4095: data <= 'd1; 4096: data <= 'd1; 4097: data <= 'd0; 4098: data <= 'd0; 4099: data <= 'd0; 4100: data <= 'd0; 4101: data <= 'd0; 4102: data <= 'd0; 4103: data <= 'd0; 4104: data <= 'd0; 4105: data <= 'd0; 4106: data <= 'd0; 4107: data <= 'd0; 4108: data <= 'd0; 4109: data <= 'd1; 4110: data <= 'd1; 4111: data <= 'd1; 4112: data <= 'd1; 4113: data <= 'd1; 4114: data <= 'd1; 4115: data <= 'd1; 4116: data <= 'd1; 4117: data <= 'd1; 4118: data <= 'd1; 4119: data <= 'd1; 4120: data <= 'd1; 4121: data <= 'd1; 4122: data <= 'd1; 4123: data <= 'd1; 4124: data <= 'd0; 4125: data <= 'd0; 4126: data <= 'd0; 4127: data <= 'd0; 4128: data <= 'd0; 4129: data <= 'd0; 4130: data <= 'd0; 4131: data <= 'd0; 4132: data <= 'd0; 4133: data <= 'd0; 4134: data <= 'd0; 4135: data <= 'd0; 4136: data <= 'd0; 4137: data <= 'd0; 4138: data <= 'd0; 4139: data <= 'd0; 4140: data <= 'd0; 4141: data <= 'd0; 4142: data <= 'd0; 4143: data <= 'd0; 4144: data <= 'd0; 4145: data <= 'd0; 4146: data <= 'd0; 4147: data <= 'd0; 4148: data <= 'd0; 4149: data <= 'd0; 4150: data <= 'd0; 4151: data <= 'd0; 4152: data <= 'd0; 4153: data <= 'd0; 4154: data <= 'd0; 4155: data <= 'd0; 4156: data <= 'd1; 4157: data <= 'd1; 4158: data <= 'd1; 4159: data <= 'd1; 4160: data <= 'd1; 4161: data <= 'd1; 4162: data <= 'd1; 4163: data <= 'd1; 4164: data <= 'd1; 4165: data <= 'd1; 4166: data <= 'd1; 4167: data <= 'd1; 4168: data <= 'd1; 4169: data <= 'd1; 4170: data <= 'd1; 4171: data <= 'd1; 4172: data <= 'd1; 4173: data <= 'd1; 4174: data <= 'd0; 4175: data <= 'd0; 4176: data <= 'd0; 4177: data <= 'd0; 4178: data <= 'd0; 4179: data <= 'd0; 4180: data <= 'd0; 4181: data <= 'd0; 4182: data <= 'd0; 4183: data <= 'd0; 4184: data <= 'd0; 4185: data <= 'd0; 4186: data <= 'd0; 4187: data <= 'd0; 4188: data <= 'd0; 4189: data <= 'd0; 4190: data <= 'd0; 4191: data <= 'd0; 4192: data <= 'd0; 4193: data <= 'd0; 4194: data <= 'd0; 4195: data <= 'd0; 4196: data <= 'd0; 4197: data <= 'd0; 4198: data <= 'd0; 4199: data <= 'd0; 4200: data <= 'd0; 4201: data <= 'd0; 4202: data <= 'd1; 4203: data <= 'd1; 4204: data <= 'd1; 4205: data <= 'd1; 4206: data <= 'd1; 4207: data <= 'd1; 4208: data <= 'd1; 4209: data <= 'd1; 4210: data <= 'd1; 4211: data <= 'd1; 4212: data <= 'd1; 4213: data <= 'd1; 4214: data <= 'd1; 4215: data <= 'd1; 4216: data <= 'd1; 4217: data <= 'd1; 4218: data <= 'd1; 4219: data <= 'd1; 4220: data <= 'd1; 4221: data <= 'd1; 4222: data <= 'd1; 4223: data <= 'd1; 4224: data <= 'd0; 4225: data <= 'd0; 4226: data <= 'd0; 4227: data <= 'd0; 4228: data <= 'd0; 4229: data <= 'd0; 4230: data <= 'd0; 4231: data <= 'd0; 4232: data <= 'd0; 4233: data <= 'd0; 4234: data <= 'd0; 4235: data <= 'd0; 4236: data <= 'd0; 4237: data <= 'd1; 4238: data <= 'd1; 4239: data <= 'd1; 4240: data <= 'd1; 4241: data <= 'd1; 4242: data <= 'd1; 4243: data <= 'd1; 4244: data <= 'd1; 4245: data <= 'd1; 4246: data <= 'd1; 4247: data <= 'd1; 4248: data <= 'd1; 4249: data <= 'd1; 4250: data <= 'd1; 4251: data <= 'd0; 4252: data <= 'd0; 4253: data <= 'd0; 4254: data <= 'd0; 4255: data <= 'd0; 4256: data <= 'd0; 4257: data <= 'd0; 4258: data <= 'd0; 4259: data <= 'd0; 4260: data <= 'd0; 4261: data <= 'd0; 4262: data <= 'd0; 4263: data <= 'd0; 4264: data <= 'd0; 4265: data <= 'd0; 4266: data <= 'd0; 4267: data <= 'd0; 4268: data <= 'd0; 4269: data <= 'd0; 4270: data <= 'd0; 4271: data <= 'd0; 4272: data <= 'd0; 4273: data <= 'd0; 4274: data <= 'd0; 4275: data <= 'd0; 4276: data <= 'd0; 4277: data <= 'd0; 4278: data <= 'd0; 4279: data <= 'd0; 4280: data <= 'd0; 4281: data <= 'd0; 4282: data <= 'd0; 4283: data <= 'd0; 4284: data <= 'd0; 4285: data <= 'd1; 4286: data <= 'd1; 4287: data <= 'd1; 4288: data <= 'd1; 4289: data <= 'd1; 4290: data <= 'd1; 4291: data <= 'd1; 4292: data <= 'd1; 4293: data <= 'd1; 4294: data <= 'd1; 4295: data <= 'd1; 4296: data <= 'd1; 4297: data <= 'd1; 4298: data <= 'd1; 4299: data <= 'd0; 4300: data <= 'd0; 4301: data <= 'd0; 4302: data <= 'd0; 4303: data <= 'd0; 4304: data <= 'd0; 4305: data <= 'd0; 4306: data <= 'd0; 4307: data <= 'd0; 4308: data <= 'd0; 4309: data <= 'd0; 4310: data <= 'd0; 4311: data <= 'd0; 4312: data <= 'd0; 4313: data <= 'd0; 4314: data <= 'd0; 4315: data <= 'd0; 4316: data <= 'd0; 4317: data <= 'd0; 4318: data <= 'd0; 4319: data <= 'd0; 4320: data <= 'd0; 4321: data <= 'd0; 4322: data <= 'd0; 4323: data <= 'd0; 4324: data <= 'd0; 4325: data <= 'd0; 4326: data <= 'd0; 4327: data <= 'd0; 4328: data <= 'd0; 4329: data <= 'd0; 4330: data <= 'd0; 4331: data <= 'd1; 4332: data <= 'd1; 4333: data <= 'd1; 4334: data <= 'd1; 4335: data <= 'd1; 4336: data <= 'd1; 4337: data <= 'd1; 4338: data <= 'd1; 4339: data <= 'd1; 4340: data <= 'd1; 4341: data <= 'd1; 4342: data <= 'd1; 4343: data <= 'd1; 4344: data <= 'd1; 4345: data <= 'd1; 4346: data <= 'd1; 4347: data <= 'd1; 4348: data <= 'd1; 4349: data <= 'd1; 4350: data <= 'd1; 4351: data <= 'd1; 4352: data <= 'd0; 4353: data <= 'd0; 4354: data <= 'd0; 4355: data <= 'd0; 4356: data <= 'd0; 4357: data <= 'd0; 4358: data <= 'd0; 4359: data <= 'd0; 4360: data <= 'd0; 4361: data <= 'd0; 4362: data <= 'd0; 4363: data <= 'd0; 4364: data <= 'd0; 4365: data <= 'd0; 4366: data <= 'd1; 4367: data <= 'd1; 4368: data <= 'd1; 4369: data <= 'd1; 4370: data <= 'd1; 4371: data <= 'd1; 4372: data <= 'd1; 4373: data <= 'd1; 4374: data <= 'd1; 4375: data <= 'd1; 4376: data <= 'd1; 4377: data <= 'd0; 4378: data <= 'd0; 4379: data <= 'd0; 4380: data <= 'd0; 4381: data <= 'd0; 4382: data <= 'd0; 4383: data <= 'd0; 4384: data <= 'd0; 4385: data <= 'd0; 4386: data <= 'd0; 4387: data <= 'd0; 4388: data <= 'd0; 4389: data <= 'd0; 4390: data <= 'd0; 4391: data <= 'd0; 4392: data <= 'd0; 4393: data <= 'd0; 4394: data <= 'd0; 4395: data <= 'd0; 4396: data <= 'd0; 4397: data <= 'd0; 4398: data <= 'd0; 4399: data <= 'd0; 4400: data <= 'd0; 4401: data <= 'd0; 4402: data <= 'd0; 4403: data <= 'd0; 4404: data <= 'd0; 4405: data <= 'd0; 4406: data <= 'd0; 4407: data <= 'd0; 4408: data <= 'd0; 4409: data <= 'd0; 4410: data <= 'd0; 4411: data <= 'd0; 4412: data <= 'd0; 4413: data <= 'd1; 4414: data <= 'd1; 4415: data <= 'd1; 4416: data <= 'd1; 4417: data <= 'd1; 4418: data <= 'd1; 4419: data <= 'd1; 4420: data <= 'd1; 4421: data <= 'd1; 4422: data <= 'd1; 4423: data <= 'd1; 4424: data <= 'd1; 4425: data <= 'd1; 4426: data <= 'd0; 4427: data <= 'd0; 4428: data <= 'd0; 4429: data <= 'd0; 4430: data <= 'd0; 4431: data <= 'd0; 4432: data <= 'd0; 4433: data <= 'd0; 4434: data <= 'd0; 4435: data <= 'd0; 4436: data <= 'd0; 4437: data <= 'd0; 4438: data <= 'd0; 4439: data <= 'd0; 4440: data <= 'd0; 4441: data <= 'd0; 4442: data <= 'd0; 4443: data <= 'd0; 4444: data <= 'd0; 4445: data <= 'd0; 4446: data <= 'd0; 4447: data <= 'd0; 4448: data <= 'd0; 4449: data <= 'd0; 4450: data <= 'd0; 4451: data <= 'd0; 4452: data <= 'd0; 4453: data <= 'd0; 4454: data <= 'd0; 4455: data <= 'd0; 4456: data <= 'd0; 4457: data <= 'd0; 4458: data <= 'd0; 4459: data <= 'd0; 4460: data <= 'd1; 4461: data <= 'd1; 4462: data <= 'd1; 4463: data <= 'd1; 4464: data <= 'd1; 4465: data <= 'd1; 4466: data <= 'd1; 4467: data <= 'd1; 4468: data <= 'd1; 4469: data <= 'd1; 4470: data <= 'd1; 4471: data <= 'd1; 4472: data <= 'd1; 4473: data <= 'd1; 4474: data <= 'd1; 4475: data <= 'd1; 4476: data <= 'd1; 4477: data <= 'd1; 4478: data <= 'd1; 4479: data <= 'd1; 4480: data <= 'd0; 4481: data <= 'd0; 4482: data <= 'd0; 4483: data <= 'd0; 4484: data <= 'd0; 4485: data <= 'd0; 4486: data <= 'd0; 4487: data <= 'd0; 4488: data <= 'd0; 4489: data <= 'd0; 4490: data <= 'd0; 4491: data <= 'd0; 4492: data <= 'd0; 4493: data <= 'd0; 4494: data <= 'd1; 4495: data <= 'd1; 4496: data <= 'd1; 4497: data <= 'd1; 4498: data <= 'd1; 4499: data <= 'd1; 4500: data <= 'd1; 4501: data <= 'd1; 4502: data <= 'd1; 4503: data <= 'd1; 4504: data <= 'd0; 4505: data <= 'd0; 4506: data <= 'd0; 4507: data <= 'd0; 4508: data <= 'd0; 4509: data <= 'd0; 4510: data <= 'd0; 4511: data <= 'd0; 4512: data <= 'd0; 4513: data <= 'd0; 4514: data <= 'd0; 4515: data <= 'd0; 4516: data <= 'd0; 4517: data <= 'd0; 4518: data <= 'd0; 4519: data <= 'd0; 4520: data <= 'd0; 4521: data <= 'd0; 4522: data <= 'd0; 4523: data <= 'd0; 4524: data <= 'd0; 4525: data <= 'd0; 4526: data <= 'd0; 4527: data <= 'd0; 4528: data <= 'd0; 4529: data <= 'd0; 4530: data <= 'd0; 4531: data <= 'd0; 4532: data <= 'd0; 4533: data <= 'd0; 4534: data <= 'd0; 4535: data <= 'd0; 4536: data <= 'd0; 4537: data <= 'd0; 4538: data <= 'd0; 4539: data <= 'd0; 4540: data <= 'd0; 4541: data <= 'd0; 4542: data <= 'd1; 4543: data <= 'd1; 4544: data <= 'd1; 4545: data <= 'd1; 4546: data <= 'd1; 4547: data <= 'd1; 4548: data <= 'd1; 4549: data <= 'd1; 4550: data <= 'd1; 4551: data <= 'd1; 4552: data <= 'd1; 4553: data <= 'd0; 4554: data <= 'd0; 4555: data <= 'd0; 4556: data <= 'd0; 4557: data <= 'd0; 4558: data <= 'd0; 4559: data <= 'd0; 4560: data <= 'd0; 4561: data <= 'd0; 4562: data <= 'd0; 4563: data <= 'd0; 4564: data <= 'd0; 4565: data <= 'd0; 4566: data <= 'd0; 4567: data <= 'd0; 4568: data <= 'd0; 4569: data <= 'd0; 4570: data <= 'd0; 4571: data <= 'd0; 4572: data <= 'd0; 4573: data <= 'd0; 4574: data <= 'd0; 4575: data <= 'd0; 4576: data <= 'd0; 4577: data <= 'd0; 4578: data <= 'd0; 4579: data <= 'd0; 4580: data <= 'd0; 4581: data <= 'd0; 4582: data <= 'd0; 4583: data <= 'd0; 4584: data <= 'd0; 4585: data <= 'd0; 4586: data <= 'd0; 4587: data <= 'd0; 4588: data <= 'd0; 4589: data <= 'd0; 4590: data <= 'd1; 4591: data <= 'd1; 4592: data <= 'd1; 4593: data <= 'd1; 4594: data <= 'd1; 4595: data <= 'd0; 4596: data <= 'd0; 4597: data <= 'd0; 4598: data <= 'd1; 4599: data <= 'd1; 4600: data <= 'd1; 4601: data <= 'd1; 4602: data <= 'd1; 4603: data <= 'd1; 4604: data <= 'd1; 4605: data <= 'd1; 4606: data <= 'd1; 4607: data <= 'd1; 4608: data <= 'd0; 4609: data <= 'd0; 4610: data <= 'd0; 4611: data <= 'd0; 4612: data <= 'd0; 4613: data <= 'd0; 4614: data <= 'd0; 4615: data <= 'd0; 4616: data <= 'd0; 4617: data <= 'd0; 4618: data <= 'd0; 4619: data <= 'd0; 4620: data <= 'd0; 4621: data <= 'd0; 4622: data <= 'd1; 4623: data <= 'd1; 4624: data <= 'd1; 4625: data <= 'd1; 4626: data <= 'd1; 4627: data <= 'd1; 4628: data <= 'd1; 4629: data <= 'd1; 4630: data <= 'd1; 4631: data <= 'd1; 4632: data <= 'd0; 4633: data <= 'd0; 4634: data <= 'd0; 4635: data <= 'd0; 4636: data <= 'd0; 4637: data <= 'd0; 4638: data <= 'd0; 4639: data <= 'd0; 4640: data <= 'd0; 4641: data <= 'd0; 4642: data <= 'd0; 4643: data <= 'd0; 4644: data <= 'd0; 4645: data <= 'd0; 4646: data <= 'd0; 4647: data <= 'd0; 4648: data <= 'd0; 4649: data <= 'd0; 4650: data <= 'd0; 4651: data <= 'd0; 4652: data <= 'd0; 4653: data <= 'd0; 4654: data <= 'd0; 4655: data <= 'd0; 4656: data <= 'd0; 4657: data <= 'd0; 4658: data <= 'd0; 4659: data <= 'd0; 4660: data <= 'd0; 4661: data <= 'd0; 4662: data <= 'd0; 4663: data <= 'd0; 4664: data <= 'd0; 4665: data <= 'd0; 4666: data <= 'd0; 4667: data <= 'd0; 4668: data <= 'd0; 4669: data <= 'd0; 4670: data <= 'd1; 4671: data <= 'd1; 4672: data <= 'd1; 4673: data <= 'd1; 4674: data <= 'd1; 4675: data <= 'd1; 4676: data <= 'd1; 4677: data <= 'd1; 4678: data <= 'd1; 4679: data <= 'd1; 4680: data <= 'd0; 4681: data <= 'd0; 4682: data <= 'd0; 4683: data <= 'd0; 4684: data <= 'd0; 4685: data <= 'd0; 4686: data <= 'd0; 4687: data <= 'd0; 4688: data <= 'd0; 4689: data <= 'd0; 4690: data <= 'd0; 4691: data <= 'd0; 4692: data <= 'd0; 4693: data <= 'd0; 4694: data <= 'd0; 4695: data <= 'd0; 4696: data <= 'd0; 4697: data <= 'd0; 4698: data <= 'd0; 4699: data <= 'd0; 4700: data <= 'd0; 4701: data <= 'd0; 4702: data <= 'd0; 4703: data <= 'd0; 4704: data <= 'd0; 4705: data <= 'd0; 4706: data <= 'd0; 4707: data <= 'd0; 4708: data <= 'd0; 4709: data <= 'd0; 4710: data <= 'd0; 4711: data <= 'd0; 4712: data <= 'd0; 4713: data <= 'd0; 4714: data <= 'd0; 4715: data <= 'd0; 4716: data <= 'd0; 4717: data <= 'd0; 4718: data <= 'd0; 4719: data <= 'd0; 4720: data <= 'd0; 4721: data <= 'd0; 4722: data <= 'd0; 4723: data <= 'd0; 4724: data <= 'd0; 4725: data <= 'd0; 4726: data <= 'd0; 4727: data <= 'd0; 4728: data <= 'd1; 4729: data <= 'd1; 4730: data <= 'd1; 4731: data <= 'd1; 4732: data <= 'd1; 4733: data <= 'd1; 4734: data <= 'd1; 4735: data <= 'd1; 4736: data <= 'd0; 4737: data <= 'd0; 4738: data <= 'd0; 4739: data <= 'd0; 4740: data <= 'd0; 4741: data <= 'd0; 4742: data <= 'd0; 4743: data <= 'd0; 4744: data <= 'd0; 4745: data <= 'd0; 4746: data <= 'd0; 4747: data <= 'd0; 4748: data <= 'd0; 4749: data <= 'd0; 4750: data <= 'd1; 4751: data <= 'd1; 4752: data <= 'd1; 4753: data <= 'd1; 4754: data <= 'd1; 4755: data <= 'd1; 4756: data <= 'd1; 4757: data <= 'd1; 4758: data <= 'd1; 4759: data <= 'd1; 4760: data <= 'd0; 4761: data <= 'd0; 4762: data <= 'd0; 4763: data <= 'd0; 4764: data <= 'd0; 4765: data <= 'd0; 4766: data <= 'd0; 4767: data <= 'd0; 4768: data <= 'd0; 4769: data <= 'd0; 4770: data <= 'd0; 4771: data <= 'd0; 4772: data <= 'd0; 4773: data <= 'd0; 4774: data <= 'd0; 4775: data <= 'd0; 4776: data <= 'd0; 4777: data <= 'd0; 4778: data <= 'd0; 4779: data <= 'd0; 4780: data <= 'd0; 4781: data <= 'd0; 4782: data <= 'd0; 4783: data <= 'd0; 4784: data <= 'd0; 4785: data <= 'd0; 4786: data <= 'd0; 4787: data <= 'd0; 4788: data <= 'd0; 4789: data <= 'd0; 4790: data <= 'd0; 4791: data <= 'd0; 4792: data <= 'd0; 4793: data <= 'd0; 4794: data <= 'd0; 4795: data <= 'd0; 4796: data <= 'd0; 4797: data <= 'd1; 4798: data <= 'd1; 4799: data <= 'd1; 4800: data <= 'd1; 4801: data <= 'd1; 4802: data <= 'd1; 4803: data <= 'd1; 4804: data <= 'd1; 4805: data <= 'd1; 4806: data <= 'd1; 4807: data <= 'd0; 4808: data <= 'd0; 4809: data <= 'd0; 4810: data <= 'd0; 4811: data <= 'd0; 4812: data <= 'd0; 4813: data <= 'd0; 4814: data <= 'd0; 4815: data <= 'd0; 4816: data <= 'd0; 4817: data <= 'd0; 4818: data <= 'd0; 4819: data <= 'd0; 4820: data <= 'd0; 4821: data <= 'd0; 4822: data <= 'd0; 4823: data <= 'd0; 4824: data <= 'd0; 4825: data <= 'd0; 4826: data <= 'd0; 4827: data <= 'd0; 4828: data <= 'd0; 4829: data <= 'd0; 4830: data <= 'd0; 4831: data <= 'd0; 4832: data <= 'd0; 4833: data <= 'd0; 4834: data <= 'd0; 4835: data <= 'd0; 4836: data <= 'd0; 4837: data <= 'd0; 4838: data <= 'd0; 4839: data <= 'd0; 4840: data <= 'd0; 4841: data <= 'd0; 4842: data <= 'd0; 4843: data <= 'd0; 4844: data <= 'd0; 4845: data <= 'd0; 4846: data <= 'd0; 4847: data <= 'd0; 4848: data <= 'd0; 4849: data <= 'd0; 4850: data <= 'd0; 4851: data <= 'd0; 4852: data <= 'd0; 4853: data <= 'd0; 4854: data <= 'd0; 4855: data <= 'd0; 4856: data <= 'd0; 4857: data <= 'd0; 4858: data <= 'd0; 4859: data <= 'd1; 4860: data <= 'd1; 4861: data <= 'd1; 4862: data <= 'd1; 4863: data <= 'd1; 4864: data <= 'd0; 4865: data <= 'd0; 4866: data <= 'd0; 4867: data <= 'd0; 4868: data <= 'd0; 4869: data <= 'd0; 4870: data <= 'd0; 4871: data <= 'd0; 4872: data <= 'd0; 4873: data <= 'd0; 4874: data <= 'd0; 4875: data <= 'd0; 4876: data <= 'd0; 4877: data <= 'd0; 4878: data <= 'd1; 4879: data <= 'd1; 4880: data <= 'd1; 4881: data <= 'd1; 4882: data <= 'd1; 4883: data <= 'd1; 4884: data <= 'd1; 4885: data <= 'd1; 4886: data <= 'd1; 4887: data <= 'd1; 4888: data <= 'd0; 4889: data <= 'd0; 4890: data <= 'd0; 4891: data <= 'd0; 4892: data <= 'd0; 4893: data <= 'd0; 4894: data <= 'd0; 4895: data <= 'd0; 4896: data <= 'd0; 4897: data <= 'd0; 4898: data <= 'd0; 4899: data <= 'd0; 4900: data <= 'd0; 4901: data <= 'd0; 4902: data <= 'd0; 4903: data <= 'd0; 4904: data <= 'd0; 4905: data <= 'd0; 4906: data <= 'd1; 4907: data <= 'd1; 4908: data <= 'd1; 4909: data <= 'd1; 4910: data <= 'd0; 4911: data <= 'd0; 4912: data <= 'd0; 4913: data <= 'd0; 4914: data <= 'd0; 4915: data <= 'd0; 4916: data <= 'd0; 4917: data <= 'd0; 4918: data <= 'd0; 4919: data <= 'd0; 4920: data <= 'd0; 4921: data <= 'd0; 4922: data <= 'd0; 4923: data <= 'd0; 4924: data <= 'd1; 4925: data <= 'd1; 4926: data <= 'd1; 4927: data <= 'd1; 4928: data <= 'd1; 4929: data <= 'd1; 4930: data <= 'd1; 4931: data <= 'd1; 4932: data <= 'd1; 4933: data <= 'd1; 4934: data <= 'd0; 4935: data <= 'd0; 4936: data <= 'd0; 4937: data <= 'd0; 4938: data <= 'd0; 4939: data <= 'd0; 4940: data <= 'd0; 4941: data <= 'd0; 4942: data <= 'd0; 4943: data <= 'd0; 4944: data <= 'd0; 4945: data <= 'd0; 4946: data <= 'd0; 4947: data <= 'd0; 4948: data <= 'd0; 4949: data <= 'd0; 4950: data <= 'd0; 4951: data <= 'd0; 4952: data <= 'd0; 4953: data <= 'd0; 4954: data <= 'd0; 4955: data <= 'd0; 4956: data <= 'd0; 4957: data <= 'd0; 4958: data <= 'd0; 4959: data <= 'd0; 4960: data <= 'd0; 4961: data <= 'd0; 4962: data <= 'd0; 4963: data <= 'd0; 4964: data <= 'd0; 4965: data <= 'd0; 4966: data <= 'd0; 4967: data <= 'd0; 4968: data <= 'd0; 4969: data <= 'd0; 4970: data <= 'd0; 4971: data <= 'd0; 4972: data <= 'd0; 4973: data <= 'd0; 4974: data <= 'd0; 4975: data <= 'd0; 4976: data <= 'd0; 4977: data <= 'd0; 4978: data <= 'd0; 4979: data <= 'd0; 4980: data <= 'd0; 4981: data <= 'd0; 4982: data <= 'd0; 4983: data <= 'd0; 4984: data <= 'd0; 4985: data <= 'd0; 4986: data <= 'd0; 4987: data <= 'd1; 4988: data <= 'd1; 4989: data <= 'd1; 4990: data <= 'd1; 4991: data <= 'd1; 4992: data <= 'd0; 4993: data <= 'd0; 4994: data <= 'd0; 4995: data <= 'd0; 4996: data <= 'd0; 4997: data <= 'd0; 4998: data <= 'd0; 4999: data <= 'd0; 5000: data <= 'd0; 5001: data <= 'd0; 5002: data <= 'd0; 5003: data <= 'd0; 5004: data <= 'd0; 5005: data <= 'd0; 5006: data <= 'd1; 5007: data <= 'd1; 5008: data <= 'd1; 5009: data <= 'd1; 5010: data <= 'd1; 5011: data <= 'd1; 5012: data <= 'd1; 5013: data <= 'd1; 5014: data <= 'd1; 5015: data <= 'd0; 5016: data <= 'd0; 5017: data <= 'd0; 5018: data <= 'd0; 5019: data <= 'd0; 5020: data <= 'd0; 5021: data <= 'd0; 5022: data <= 'd0; 5023: data <= 'd0; 5024: data <= 'd0; 5025: data <= 'd0; 5026: data <= 'd0; 5027: data <= 'd0; 5028: data <= 'd0; 5029: data <= 'd0; 5030: data <= 'd0; 5031: data <= 'd0; 5032: data <= 'd0; 5033: data <= 'd0; 5034: data <= 'd0; 5035: data <= 'd0; 5036: data <= 'd0; 5037: data <= 'd1; 5038: data <= 'd1; 5039: data <= 'd0; 5040: data <= 'd0; 5041: data <= 'd1; 5042: data <= 'd1; 5043: data <= 'd1; 5044: data <= 'd1; 5045: data <= 'd0; 5046: data <= 'd0; 5047: data <= 'd0; 5048: data <= 'd0; 5049: data <= 'd0; 5050: data <= 'd1; 5051: data <= 'd1; 5052: data <= 'd1; 5053: data <= 'd1; 5054: data <= 'd1; 5055: data <= 'd1; 5056: data <= 'd1; 5057: data <= 'd1; 5058: data <= 'd1; 5059: data <= 'd1; 5060: data <= 'd1; 5061: data <= 'd0; 5062: data <= 'd0; 5063: data <= 'd0; 5064: data <= 'd0; 5065: data <= 'd0; 5066: data <= 'd0; 5067: data <= 'd0; 5068: data <= 'd0; 5069: data <= 'd0; 5070: data <= 'd0; 5071: data <= 'd0; 5072: data <= 'd0; 5073: data <= 'd0; 5074: data <= 'd0; 5075: data <= 'd0; 5076: data <= 'd0; 5077: data <= 'd0; 5078: data <= 'd0; 5079: data <= 'd0; 5080: data <= 'd0; 5081: data <= 'd0; 5082: data <= 'd0; 5083: data <= 'd0; 5084: data <= 'd0; 5085: data <= 'd0; 5086: data <= 'd0; 5087: data <= 'd0; 5088: data <= 'd0; 5089: data <= 'd0; 5090: data <= 'd0; 5091: data <= 'd0; 5092: data <= 'd0; 5093: data <= 'd0; 5094: data <= 'd0; 5095: data <= 'd0; 5096: data <= 'd0; 5097: data <= 'd0; 5098: data <= 'd0; 5099: data <= 'd0; 5100: data <= 'd0; 5101: data <= 'd0; 5102: data <= 'd0; 5103: data <= 'd0; 5104: data <= 'd0; 5105: data <= 'd0; 5106: data <= 'd0; 5107: data <= 'd0; 5108: data <= 'd0; 5109: data <= 'd0; 5110: data <= 'd0; 5111: data <= 'd0; 5112: data <= 'd0; 5113: data <= 'd0; 5114: data <= 'd0; 5115: data <= 'd1; 5116: data <= 'd1; 5117: data <= 'd1; 5118: data <= 'd1; 5119: data <= 'd1; 5120: data <= 'd0; 5121: data <= 'd0; 5122: data <= 'd0; 5123: data <= 'd0; 5124: data <= 'd0; 5125: data <= 'd0; 5126: data <= 'd0; 5127: data <= 'd0; 5128: data <= 'd0; 5129: data <= 'd0; 5130: data <= 'd0; 5131: data <= 'd0; 5132: data <= 'd0; 5133: data <= 'd0; 5134: data <= 'd1; 5135: data <= 'd1; 5136: data <= 'd1; 5137: data <= 'd1; 5138: data <= 'd1; 5139: data <= 'd1; 5140: data <= 'd1; 5141: data <= 'd1; 5142: data <= 'd1; 5143: data <= 'd0; 5144: data <= 'd0; 5145: data <= 'd0; 5146: data <= 'd0; 5147: data <= 'd0; 5148: data <= 'd0; 5149: data <= 'd0; 5150: data <= 'd0; 5151: data <= 'd0; 5152: data <= 'd0; 5153: data <= 'd0; 5154: data <= 'd0; 5155: data <= 'd0; 5156: data <= 'd0; 5157: data <= 'd0; 5158: data <= 'd0; 5159: data <= 'd0; 5160: data <= 'd0; 5161: data <= 'd0; 5162: data <= 'd0; 5163: data <= 'd0; 5164: data <= 'd0; 5165: data <= 'd0; 5166: data <= 'd1; 5167: data <= 'd1; 5168: data <= 'd1; 5169: data <= 'd1; 5170: data <= 'd1; 5171: data <= 'd1; 5172: data <= 'd1; 5173: data <= 'd1; 5174: data <= 'd1; 5175: data <= 'd1; 5176: data <= 'd1; 5177: data <= 'd1; 5178: data <= 'd1; 5179: data <= 'd1; 5180: data <= 'd1; 5181: data <= 'd1; 5182: data <= 'd1; 5183: data <= 'd1; 5184: data <= 'd1; 5185: data <= 'd1; 5186: data <= 'd1; 5187: data <= 'd1; 5188: data <= 'd0; 5189: data <= 'd0; 5190: data <= 'd0; 5191: data <= 'd0; 5192: data <= 'd0; 5193: data <= 'd0; 5194: data <= 'd0; 5195: data <= 'd0; 5196: data <= 'd0; 5197: data <= 'd0; 5198: data <= 'd0; 5199: data <= 'd0; 5200: data <= 'd0; 5201: data <= 'd0; 5202: data <= 'd0; 5203: data <= 'd0; 5204: data <= 'd0; 5205: data <= 'd0; 5206: data <= 'd0; 5207: data <= 'd0; 5208: data <= 'd0; 5209: data <= 'd0; 5210: data <= 'd0; 5211: data <= 'd0; 5212: data <= 'd0; 5213: data <= 'd0; 5214: data <= 'd0; 5215: data <= 'd0; 5216: data <= 'd0; 5217: data <= 'd0; 5218: data <= 'd0; 5219: data <= 'd0; 5220: data <= 'd0; 5221: data <= 'd0; 5222: data <= 'd0; 5223: data <= 'd0; 5224: data <= 'd0; 5225: data <= 'd0; 5226: data <= 'd0; 5227: data <= 'd0; 5228: data <= 'd0; 5229: data <= 'd0; 5230: data <= 'd0; 5231: data <= 'd0; 5232: data <= 'd0; 5233: data <= 'd0; 5234: data <= 'd0; 5235: data <= 'd0; 5236: data <= 'd0; 5237: data <= 'd0; 5238: data <= 'd0; 5239: data <= 'd0; 5240: data <= 'd0; 5241: data <= 'd0; 5242: data <= 'd0; 5243: data <= 'd0; 5244: data <= 'd1; 5245: data <= 'd1; 5246: data <= 'd1; 5247: data <= 'd1; 5248: data <= 'd0; 5249: data <= 'd0; 5250: data <= 'd0; 5251: data <= 'd0; 5252: data <= 'd0; 5253: data <= 'd0; 5254: data <= 'd0; 5255: data <= 'd0; 5256: data <= 'd0; 5257: data <= 'd0; 5258: data <= 'd0; 5259: data <= 'd0; 5260: data <= 'd0; 5261: data <= 'd0; 5262: data <= 'd1; 5263: data <= 'd1; 5264: data <= 'd1; 5265: data <= 'd1; 5266: data <= 'd1; 5267: data <= 'd1; 5268: data <= 'd1; 5269: data <= 'd1; 5270: data <= 'd1; 5271: data <= 'd0; 5272: data <= 'd0; 5273: data <= 'd0; 5274: data <= 'd0; 5275: data <= 'd0; 5276: data <= 'd0; 5277: data <= 'd0; 5278: data <= 'd0; 5279: data <= 'd0; 5280: data <= 'd0; 5281: data <= 'd0; 5282: data <= 'd0; 5283: data <= 'd0; 5284: data <= 'd0; 5285: data <= 'd0; 5286: data <= 'd0; 5287: data <= 'd0; 5288: data <= 'd0; 5289: data <= 'd0; 5290: data <= 'd0; 5291: data <= 'd0; 5292: data <= 'd0; 5293: data <= 'd0; 5294: data <= 'd0; 5295: data <= 'd1; 5296: data <= 'd1; 5297: data <= 'd1; 5298: data <= 'd1; 5299: data <= 'd1; 5300: data <= 'd1; 5301: data <= 'd1; 5302: data <= 'd1; 5303: data <= 'd1; 5304: data <= 'd1; 5305: data <= 'd1; 5306: data <= 'd1; 5307: data <= 'd1; 5308: data <= 'd1; 5309: data <= 'd1; 5310: data <= 'd1; 5311: data <= 'd1; 5312: data <= 'd1; 5313: data <= 'd1; 5314: data <= 'd1; 5315: data <= 'd0; 5316: data <= 'd0; 5317: data <= 'd0; 5318: data <= 'd0; 5319: data <= 'd0; 5320: data <= 'd0; 5321: data <= 'd0; 5322: data <= 'd0; 5323: data <= 'd0; 5324: data <= 'd0; 5325: data <= 'd0; 5326: data <= 'd0; 5327: data <= 'd0; 5328: data <= 'd0; 5329: data <= 'd0; 5330: data <= 'd0; 5331: data <= 'd0; 5332: data <= 'd0; 5333: data <= 'd0; 5334: data <= 'd0; 5335: data <= 'd0; 5336: data <= 'd0; 5337: data <= 'd0; 5338: data <= 'd0; 5339: data <= 'd0; 5340: data <= 'd0; 5341: data <= 'd0; 5342: data <= 'd0; 5343: data <= 'd0; 5344: data <= 'd0; 5345: data <= 'd0; 5346: data <= 'd0; 5347: data <= 'd0; 5348: data <= 'd0; 5349: data <= 'd0; 5350: data <= 'd0; 5351: data <= 'd0; 5352: data <= 'd0; 5353: data <= 'd0; 5354: data <= 'd0; 5355: data <= 'd0; 5356: data <= 'd0; 5357: data <= 'd0; 5358: data <= 'd0; 5359: data <= 'd0; 5360: data <= 'd0; 5361: data <= 'd0; 5362: data <= 'd0; 5363: data <= 'd0; 5364: data <= 'd0; 5365: data <= 'd0; 5366: data <= 'd0; 5367: data <= 'd0; 5368: data <= 'd0; 5369: data <= 'd0; 5370: data <= 'd0; 5371: data <= 'd0; 5372: data <= 'd1; 5373: data <= 'd1; 5374: data <= 'd1; 5375: data <= 'd1; 5376: data <= 'd0; 5377: data <= 'd0; 5378: data <= 'd0; 5379: data <= 'd0; 5380: data <= 'd0; 5381: data <= 'd0; 5382: data <= 'd0; 5383: data <= 'd0; 5384: data <= 'd0; 5385: data <= 'd0; 5386: data <= 'd0; 5387: data <= 'd0; 5388: data <= 'd0; 5389: data <= 'd1; 5390: data <= 'd1; 5391: data <= 'd1; 5392: data <= 'd1; 5393: data <= 'd1; 5394: data <= 'd1; 5395: data <= 'd1; 5396: data <= 'd1; 5397: data <= 'd1; 5398: data <= 'd1; 5399: data <= 'd0; 5400: data <= 'd0; 5401: data <= 'd0; 5402: data <= 'd0; 5403: data <= 'd0; 5404: data <= 'd0; 5405: data <= 'd0; 5406: data <= 'd0; 5407: data <= 'd0; 5408: data <= 'd0; 5409: data <= 'd0; 5410: data <= 'd0; 5411: data <= 'd0; 5412: data <= 'd0; 5413: data <= 'd0; 5414: data <= 'd0; 5415: data <= 'd0; 5416: data <= 'd0; 5417: data <= 'd0; 5418: data <= 'd0; 5419: data <= 'd0; 5420: data <= 'd0; 5421: data <= 'd0; 5422: data <= 'd1; 5423: data <= 'd1; 5424: data <= 'd1; 5425: data <= 'd0; 5426: data <= 'd0; 5427: data <= 'd1; 5428: data <= 'd1; 5429: data <= 'd1; 5430: data <= 'd1; 5431: data <= 'd1; 5432: data <= 'd1; 5433: data <= 'd1; 5434: data <= 'd1; 5435: data <= 'd1; 5436: data <= 'd1; 5437: data <= 'd1; 5438: data <= 'd1; 5439: data <= 'd1; 5440: data <= 'd1; 5441: data <= 'd1; 5442: data <= 'd1; 5443: data <= 'd0; 5444: data <= 'd0; 5445: data <= 'd0; 5446: data <= 'd0; 5447: data <= 'd0; 5448: data <= 'd0; 5449: data <= 'd0; 5450: data <= 'd0; 5451: data <= 'd0; 5452: data <= 'd0; 5453: data <= 'd0; 5454: data <= 'd0; 5455: data <= 'd0; 5456: data <= 'd0; 5457: data <= 'd0; 5458: data <= 'd0; 5459: data <= 'd0; 5460: data <= 'd0; 5461: data <= 'd0; 5462: data <= 'd0; 5463: data <= 'd0; 5464: data <= 'd0; 5465: data <= 'd0; 5466: data <= 'd0; 5467: data <= 'd0; 5468: data <= 'd0; 5469: data <= 'd0; 5470: data <= 'd0; 5471: data <= 'd0; 5472: data <= 'd0; 5473: data <= 'd0; 5474: data <= 'd0; 5475: data <= 'd0; 5476: data <= 'd0; 5477: data <= 'd0; 5478: data <= 'd0; 5479: data <= 'd0; 5480: data <= 'd0; 5481: data <= 'd0; 5482: data <= 'd0; 5483: data <= 'd0; 5484: data <= 'd0; 5485: data <= 'd0; 5486: data <= 'd0; 5487: data <= 'd0; 5488: data <= 'd0; 5489: data <= 'd0; 5490: data <= 'd0; 5491: data <= 'd0; 5492: data <= 'd0; 5493: data <= 'd0; 5494: data <= 'd0; 5495: data <= 'd0; 5496: data <= 'd0; 5497: data <= 'd0; 5498: data <= 'd0; 5499: data <= 'd0; 5500: data <= 'd0; 5501: data <= 'd1; 5502: data <= 'd1; 5503: data <= 'd1; 5504: data <= 'd0; 5505: data <= 'd0; 5506: data <= 'd0; 5507: data <= 'd0; 5508: data <= 'd0; 5509: data <= 'd0; 5510: data <= 'd0; 5511: data <= 'd0; 5512: data <= 'd0; 5513: data <= 'd0; 5514: data <= 'd0; 5515: data <= 'd0; 5516: data <= 'd0; 5517: data <= 'd1; 5518: data <= 'd1; 5519: data <= 'd1; 5520: data <= 'd1; 5521: data <= 'd1; 5522: data <= 'd1; 5523: data <= 'd1; 5524: data <= 'd1; 5525: data <= 'd1; 5526: data <= 'd0; 5527: data <= 'd0; 5528: data <= 'd0; 5529: data <= 'd0; 5530: data <= 'd0; 5531: data <= 'd0; 5532: data <= 'd0; 5533: data <= 'd0; 5534: data <= 'd0; 5535: data <= 'd0; 5536: data <= 'd0; 5537: data <= 'd0; 5538: data <= 'd0; 5539: data <= 'd0; 5540: data <= 'd0; 5541: data <= 'd0; 5542: data <= 'd0; 5543: data <= 'd0; 5544: data <= 'd0; 5545: data <= 'd0; 5546: data <= 'd0; 5547: data <= 'd0; 5548: data <= 'd0; 5549: data <= 'd0; 5550: data <= 'd1; 5551: data <= 'd1; 5552: data <= 'd0; 5553: data <= 'd0; 5554: data <= 'd0; 5555: data <= 'd0; 5556: data <= 'd0; 5557: data <= 'd0; 5558: data <= 'd1; 5559: data <= 'd1; 5560: data <= 'd1; 5561: data <= 'd1; 5562: data <= 'd1; 5563: data <= 'd1; 5564: data <= 'd1; 5565: data <= 'd1; 5566: data <= 'd1; 5567: data <= 'd1; 5568: data <= 'd1; 5569: data <= 'd1; 5570: data <= 'd1; 5571: data <= 'd0; 5572: data <= 'd0; 5573: data <= 'd0; 5574: data <= 'd0; 5575: data <= 'd0; 5576: data <= 'd0; 5577: data <= 'd0; 5578: data <= 'd0; 5579: data <= 'd0; 5580: data <= 'd0; 5581: data <= 'd0; 5582: data <= 'd0; 5583: data <= 'd0; 5584: data <= 'd0; 5585: data <= 'd0; 5586: data <= 'd0; 5587: data <= 'd0; 5588: data <= 'd0; 5589: data <= 'd0; 5590: data <= 'd0; 5591: data <= 'd0; 5592: data <= 'd0; 5593: data <= 'd0; 5594: data <= 'd0; 5595: data <= 'd0; 5596: data <= 'd0; 5597: data <= 'd0; 5598: data <= 'd0; 5599: data <= 'd0; 5600: data <= 'd0; 5601: data <= 'd0; 5602: data <= 'd0; 5603: data <= 'd0; 5604: data <= 'd0; 5605: data <= 'd0; 5606: data <= 'd0; 5607: data <= 'd0; 5608: data <= 'd0; 5609: data <= 'd0; 5610: data <= 'd0; 5611: data <= 'd0; 5612: data <= 'd0; 5613: data <= 'd0; 5614: data <= 'd0; 5615: data <= 'd0; 5616: data <= 'd0; 5617: data <= 'd0; 5618: data <= 'd0; 5619: data <= 'd0; 5620: data <= 'd0; 5621: data <= 'd0; 5622: data <= 'd0; 5623: data <= 'd0; 5624: data <= 'd0; 5625: data <= 'd0; 5626: data <= 'd0; 5627: data <= 'd0; 5628: data <= 'd0; 5629: data <= 'd1; 5630: data <= 'd1; 5631: data <= 'd1; 5632: data <= 'd0; 5633: data <= 'd0; 5634: data <= 'd0; 5635: data <= 'd0; 5636: data <= 'd0; 5637: data <= 'd0; 5638: data <= 'd0; 5639: data <= 'd0; 5640: data <= 'd0; 5641: data <= 'd0; 5642: data <= 'd0; 5643: data <= 'd0; 5644: data <= 'd0; 5645: data <= 'd1; 5646: data <= 'd1; 5647: data <= 'd1; 5648: data <= 'd1; 5649: data <= 'd1; 5650: data <= 'd1; 5651: data <= 'd1; 5652: data <= 'd1; 5653: data <= 'd1; 5654: data <= 'd1; 5655: data <= 'd0; 5656: data <= 'd0; 5657: data <= 'd0; 5658: data <= 'd0; 5659: data <= 'd0; 5660: data <= 'd0; 5661: data <= 'd0; 5662: data <= 'd0; 5663: data <= 'd0; 5664: data <= 'd0; 5665: data <= 'd0; 5666: data <= 'd0; 5667: data <= 'd0; 5668: data <= 'd0; 5669: data <= 'd0; 5670: data <= 'd0; 5671: data <= 'd0; 5672: data <= 'd0; 5673: data <= 'd0; 5674: data <= 'd0; 5675: data <= 'd0; 5676: data <= 'd0; 5677: data <= 'd0; 5678: data <= 'd1; 5679: data <= 'd0; 5680: data <= 'd0; 5681: data <= 'd0; 5682: data <= 'd0; 5683: data <= 'd0; 5684: data <= 'd0; 5685: data <= 'd0; 5686: data <= 'd1; 5687: data <= 'd1; 5688: data <= 'd1; 5689: data <= 'd1; 5690: data <= 'd1; 5691: data <= 'd0; 5692: data <= 'd0; 5693: data <= 'd0; 5694: data <= 'd0; 5695: data <= 'd1; 5696: data <= 'd1; 5697: data <= 'd1; 5698: data <= 'd1; 5699: data <= 'd1; 5700: data <= 'd0; 5701: data <= 'd0; 5702: data <= 'd0; 5703: data <= 'd0; 5704: data <= 'd0; 5705: data <= 'd0; 5706: data <= 'd0; 5707: data <= 'd0; 5708: data <= 'd0; 5709: data <= 'd0; 5710: data <= 'd0; 5711: data <= 'd0; 5712: data <= 'd0; 5713: data <= 'd0; 5714: data <= 'd0; 5715: data <= 'd0; 5716: data <= 'd0; 5717: data <= 'd0; 5718: data <= 'd0; 5719: data <= 'd0; 5720: data <= 'd0; 5721: data <= 'd0; 5722: data <= 'd0; 5723: data <= 'd0; 5724: data <= 'd0; 5725: data <= 'd0; 5726: data <= 'd0; 5727: data <= 'd0; 5728: data <= 'd0; 5729: data <= 'd0; 5730: data <= 'd0; 5731: data <= 'd0; 5732: data <= 'd0; 5733: data <= 'd0; 5734: data <= 'd0; 5735: data <= 'd0; 5736: data <= 'd0; 5737: data <= 'd0; 5738: data <= 'd0; 5739: data <= 'd0; 5740: data <= 'd0; 5741: data <= 'd0; 5742: data <= 'd0; 5743: data <= 'd0; 5744: data <= 'd0; 5745: data <= 'd0; 5746: data <= 'd0; 5747: data <= 'd0; 5748: data <= 'd0; 5749: data <= 'd0; 5750: data <= 'd0; 5751: data <= 'd0; 5752: data <= 'd0; 5753: data <= 'd0; 5754: data <= 'd0; 5755: data <= 'd0; 5756: data <= 'd0; 5757: data <= 'd0; 5758: data <= 'd1; 5759: data <= 'd1; 5760: data <= 'd0; 5761: data <= 'd0; 5762: data <= 'd0; 5763: data <= 'd0; 5764: data <= 'd0; 5765: data <= 'd0; 5766: data <= 'd0; 5767: data <= 'd0; 5768: data <= 'd0; 5769: data <= 'd0; 5770: data <= 'd0; 5771: data <= 'd0; 5772: data <= 'd0; 5773: data <= 'd1; 5774: data <= 'd1; 5775: data <= 'd1; 5776: data <= 'd1; 5777: data <= 'd1; 5778: data <= 'd1; 5779: data <= 'd1; 5780: data <= 'd1; 5781: data <= 'd1; 5782: data <= 'd1; 5783: data <= 'd1; 5784: data <= 'd0; 5785: data <= 'd0; 5786: data <= 'd0; 5787: data <= 'd0; 5788: data <= 'd0; 5789: data <= 'd0; 5790: data <= 'd0; 5791: data <= 'd0; 5792: data <= 'd0; 5793: data <= 'd0; 5794: data <= 'd0; 5795: data <= 'd0; 5796: data <= 'd0; 5797: data <= 'd0; 5798: data <= 'd0; 5799: data <= 'd0; 5800: data <= 'd0; 5801: data <= 'd0; 5802: data <= 'd0; 5803: data <= 'd0; 5804: data <= 'd0; 5805: data <= 'd0; 5806: data <= 'd0; 5807: data <= 'd0; 5808: data <= 'd0; 5809: data <= 'd0; 5810: data <= 'd0; 5811: data <= 'd0; 5812: data <= 'd0; 5813: data <= 'd1; 5814: data <= 'd1; 5815: data <= 'd1; 5816: data <= 'd1; 5817: data <= 'd1; 5818: data <= 'd0; 5819: data <= 'd0; 5820: data <= 'd0; 5821: data <= 'd0; 5822: data <= 'd0; 5823: data <= 'd0; 5824: data <= 'd1; 5825: data <= 'd1; 5826: data <= 'd1; 5827: data <= 'd1; 5828: data <= 'd0; 5829: data <= 'd0; 5830: data <= 'd0; 5831: data <= 'd0; 5832: data <= 'd0; 5833: data <= 'd0; 5834: data <= 'd0; 5835: data <= 'd0; 5836: data <= 'd0; 5837: data <= 'd0; 5838: data <= 'd0; 5839: data <= 'd0; 5840: data <= 'd0; 5841: data <= 'd0; 5842: data <= 'd0; 5843: data <= 'd0; 5844: data <= 'd0; 5845: data <= 'd0; 5846: data <= 'd0; 5847: data <= 'd0; 5848: data <= 'd0; 5849: data <= 'd0; 5850: data <= 'd0; 5851: data <= 'd0; 5852: data <= 'd0; 5853: data <= 'd0; 5854: data <= 'd0; 5855: data <= 'd0; 5856: data <= 'd0; 5857: data <= 'd0; 5858: data <= 'd0; 5859: data <= 'd0; 5860: data <= 'd0; 5861: data <= 'd0; 5862: data <= 'd0; 5863: data <= 'd0; 5864: data <= 'd0; 5865: data <= 'd0; 5866: data <= 'd0; 5867: data <= 'd0; 5868: data <= 'd0; 5869: data <= 'd0; 5870: data <= 'd0; 5871: data <= 'd0; 5872: data <= 'd0; 5873: data <= 'd0; 5874: data <= 'd0; 5875: data <= 'd0; 5876: data <= 'd0; 5877: data <= 'd0; 5878: data <= 'd0; 5879: data <= 'd0; 5880: data <= 'd0; 5881: data <= 'd0; 5882: data <= 'd0; 5883: data <= 'd0; 5884: data <= 'd0; 5885: data <= 'd0; 5886: data <= 'd1; 5887: data <= 'd1; 5888: data <= 'd0; 5889: data <= 'd0; 5890: data <= 'd0; 5891: data <= 'd0; 5892: data <= 'd0; 5893: data <= 'd0; 5894: data <= 'd0; 5895: data <= 'd0; 5896: data <= 'd0; 5897: data <= 'd0; 5898: data <= 'd0; 5899: data <= 'd0; 5900: data <= 'd0; 5901: data <= 'd1; 5902: data <= 'd1; 5903: data <= 'd1; 5904: data <= 'd1; 5905: data <= 'd1; 5906: data <= 'd1; 5907: data <= 'd1; 5908: data <= 'd1; 5909: data <= 'd1; 5910: data <= 'd1; 5911: data <= 'd1; 5912: data <= 'd1; 5913: data <= 'd0; 5914: data <= 'd0; 5915: data <= 'd0; 5916: data <= 'd0; 5917: data <= 'd0; 5918: data <= 'd0; 5919: data <= 'd0; 5920: data <= 'd0; 5921: data <= 'd0; 5922: data <= 'd0; 5923: data <= 'd0; 5924: data <= 'd0; 5925: data <= 'd0; 5926: data <= 'd0; 5927: data <= 'd0; 5928: data <= 'd0; 5929: data <= 'd0; 5930: data <= 'd0; 5931: data <= 'd0; 5932: data <= 'd0; 5933: data <= 'd0; 5934: data <= 'd0; 5935: data <= 'd0; 5936: data <= 'd0; 5937: data <= 'd0; 5938: data <= 'd0; 5939: data <= 'd0; 5940: data <= 'd1; 5941: data <= 'd1; 5942: data <= 'd1; 5943: data <= 'd1; 5944: data <= 'd1; 5945: data <= 'd0; 5946: data <= 'd0; 5947: data <= 'd0; 5948: data <= 'd0; 5949: data <= 'd0; 5950: data <= 'd0; 5951: data <= 'd0; 5952: data <= 'd0; 5953: data <= 'd1; 5954: data <= 'd1; 5955: data <= 'd0; 5956: data <= 'd0; 5957: data <= 'd0; 5958: data <= 'd0; 5959: data <= 'd0; 5960: data <= 'd0; 5961: data <= 'd0; 5962: data <= 'd0; 5963: data <= 'd0; 5964: data <= 'd0; 5965: data <= 'd0; 5966: data <= 'd0; 5967: data <= 'd0; 5968: data <= 'd0; 5969: data <= 'd0; 5970: data <= 'd0; 5971: data <= 'd0; 5972: data <= 'd0; 5973: data <= 'd0; 5974: data <= 'd0; 5975: data <= 'd0; 5976: data <= 'd0; 5977: data <= 'd0; 5978: data <= 'd0; 5979: data <= 'd0; 5980: data <= 'd0; 5981: data <= 'd0; 5982: data <= 'd0; 5983: data <= 'd0; 5984: data <= 'd0; 5985: data <= 'd0; 5986: data <= 'd0; 5987: data <= 'd0; 5988: data <= 'd0; 5989: data <= 'd0; 5990: data <= 'd0; 5991: data <= 'd0; 5992: data <= 'd0; 5993: data <= 'd0; 5994: data <= 'd0; 5995: data <= 'd0; 5996: data <= 'd0; 5997: data <= 'd0; 5998: data <= 'd0; 5999: data <= 'd0; 6000: data <= 'd0; 6001: data <= 'd0; 6002: data <= 'd0; 6003: data <= 'd0; 6004: data <= 'd0; 6005: data <= 'd0; 6006: data <= 'd0; 6007: data <= 'd0; 6008: data <= 'd0; 6009: data <= 'd0; 6010: data <= 'd0; 6011: data <= 'd0; 6012: data <= 'd0; 6013: data <= 'd0; 6014: data <= 'd0; 6015: data <= 'd1; 6016: data <= 'd0; 6017: data <= 'd0; 6018: data <= 'd0; 6019: data <= 'd0; 6020: data <= 'd0; 6021: data <= 'd0; 6022: data <= 'd0; 6023: data <= 'd0; 6024: data <= 'd0; 6025: data <= 'd0; 6026: data <= 'd0; 6027: data <= 'd0; 6028: data <= 'd1; 6029: data <= 'd1; 6030: data <= 'd1; 6031: data <= 'd1; 6032: data <= 'd1; 6033: data <= 'd1; 6034: data <= 'd1; 6035: data <= 'd1; 6036: data <= 'd1; 6037: data <= 'd1; 6038: data <= 'd1; 6039: data <= 'd1; 6040: data <= 'd1; 6041: data <= 'd0; 6042: data <= 'd0; 6043: data <= 'd0; 6044: data <= 'd0; 6045: data <= 'd0; 6046: data <= 'd0; 6047: data <= 'd0; 6048: data <= 'd0; 6049: data <= 'd0; 6050: data <= 'd0; 6051: data <= 'd0; 6052: data <= 'd0; 6053: data <= 'd0; 6054: data <= 'd0; 6055: data <= 'd0; 6056: data <= 'd0; 6057: data <= 'd0; 6058: data <= 'd0; 6059: data <= 'd0; 6060: data <= 'd0; 6061: data <= 'd0; 6062: data <= 'd0; 6063: data <= 'd0; 6064: data <= 'd0; 6065: data <= 'd0; 6066: data <= 'd0; 6067: data <= 'd0; 6068: data <= 'd1; 6069: data <= 'd1; 6070: data <= 'd1; 6071: data <= 'd1; 6072: data <= 'd1; 6073: data <= 'd0; 6074: data <= 'd0; 6075: data <= 'd0; 6076: data <= 'd0; 6077: data <= 'd0; 6078: data <= 'd0; 6079: data <= 'd0; 6080: data <= 'd0; 6081: data <= 'd0; 6082: data <= 'd0; 6083: data <= 'd0; 6084: data <= 'd0; 6085: data <= 'd0; 6086: data <= 'd0; 6087: data <= 'd0; 6088: data <= 'd0; 6089: data <= 'd0; 6090: data <= 'd0; 6091: data <= 'd0; 6092: data <= 'd0; 6093: data <= 'd0; 6094: data <= 'd0; 6095: data <= 'd0; 6096: data <= 'd0; 6097: data <= 'd0; 6098: data <= 'd0; 6099: data <= 'd0; 6100: data <= 'd0; 6101: data <= 'd0; 6102: data <= 'd0; 6103: data <= 'd0; 6104: data <= 'd0; 6105: data <= 'd0; 6106: data <= 'd0; 6107: data <= 'd0; 6108: data <= 'd0; 6109: data <= 'd0; 6110: data <= 'd0; 6111: data <= 'd0; 6112: data <= 'd0; 6113: data <= 'd0; 6114: data <= 'd0; 6115: data <= 'd0; 6116: data <= 'd0; 6117: data <= 'd0; 6118: data <= 'd0; 6119: data <= 'd0; 6120: data <= 'd0; 6121: data <= 'd0; 6122: data <= 'd0; 6123: data <= 'd0; 6124: data <= 'd0; 6125: data <= 'd0; 6126: data <= 'd0; 6127: data <= 'd0; 6128: data <= 'd0; 6129: data <= 'd0; 6130: data <= 'd0; 6131: data <= 'd0; 6132: data <= 'd0; 6133: data <= 'd0; 6134: data <= 'd0; 6135: data <= 'd0; 6136: data <= 'd0; 6137: data <= 'd0; 6138: data <= 'd0; 6139: data <= 'd0; 6140: data <= 'd0; 6141: data <= 'd0; 6142: data <= 'd0; 6143: data <= 'd1; 6144: data <= 'd0; 6145: data <= 'd0; 6146: data <= 'd0; 6147: data <= 'd0; 6148: data <= 'd0; 6149: data <= 'd0; 6150: data <= 'd0; 6151: data <= 'd0; 6152: data <= 'd0; 6153: data <= 'd0; 6154: data <= 'd0; 6155: data <= 'd0; 6156: data <= 'd1; 6157: data <= 'd1; 6158: data <= 'd1; 6159: data <= 'd1; 6160: data <= 'd1; 6161: data <= 'd1; 6162: data <= 'd1; 6163: data <= 'd1; 6164: data <= 'd1; 6165: data <= 'd1; 6166: data <= 'd1; 6167: data <= 'd1; 6168: data <= 'd1; 6169: data <= 'd1; 6170: data <= 'd0; 6171: data <= 'd0; 6172: data <= 'd0; 6173: data <= 'd0; 6174: data <= 'd0; 6175: data <= 'd0; 6176: data <= 'd0; 6177: data <= 'd0; 6178: data <= 'd0; 6179: data <= 'd0; 6180: data <= 'd0; 6181: data <= 'd0; 6182: data <= 'd0; 6183: data <= 'd0; 6184: data <= 'd0; 6185: data <= 'd0; 6186: data <= 'd0; 6187: data <= 'd0; 6188: data <= 'd0; 6189: data <= 'd0; 6190: data <= 'd0; 6191: data <= 'd0; 6192: data <= 'd0; 6193: data <= 'd0; 6194: data <= 'd0; 6195: data <= 'd1; 6196: data <= 'd1; 6197: data <= 'd1; 6198: data <= 'd1; 6199: data <= 'd1; 6200: data <= 'd0; 6201: data <= 'd0; 6202: data <= 'd0; 6203: data <= 'd0; 6204: data <= 'd0; 6205: data <= 'd0; 6206: data <= 'd0; 6207: data <= 'd0; 6208: data <= 'd0; 6209: data <= 'd0; 6210: data <= 'd0; 6211: data <= 'd0; 6212: data <= 'd0; 6213: data <= 'd0; 6214: data <= 'd0; 6215: data <= 'd0; 6216: data <= 'd0; 6217: data <= 'd0; 6218: data <= 'd0; 6219: data <= 'd0; 6220: data <= 'd0; 6221: data <= 'd0; 6222: data <= 'd0; 6223: data <= 'd0; 6224: data <= 'd0; 6225: data <= 'd0; 6226: data <= 'd0; 6227: data <= 'd0; 6228: data <= 'd0; 6229: data <= 'd0; 6230: data <= 'd0; 6231: data <= 'd0; 6232: data <= 'd0; 6233: data <= 'd0; 6234: data <= 'd0; 6235: data <= 'd0; 6236: data <= 'd0; 6237: data <= 'd0; 6238: data <= 'd0; 6239: data <= 'd0; 6240: data <= 'd0; 6241: data <= 'd0; 6242: data <= 'd0; 6243: data <= 'd0; 6244: data <= 'd0; 6245: data <= 'd0; 6246: data <= 'd0; 6247: data <= 'd0; 6248: data <= 'd0; 6249: data <= 'd0; 6250: data <= 'd0; 6251: data <= 'd0; 6252: data <= 'd0; 6253: data <= 'd0; 6254: data <= 'd0; 6255: data <= 'd0; 6256: data <= 'd0; 6257: data <= 'd0; 6258: data <= 'd0; 6259: data <= 'd0; 6260: data <= 'd0; 6261: data <= 'd0; 6262: data <= 'd0; 6263: data <= 'd0; 6264: data <= 'd0; 6265: data <= 'd0; 6266: data <= 'd0; 6267: data <= 'd0; 6268: data <= 'd0; 6269: data <= 'd0; 6270: data <= 'd0; 6271: data <= 'd0; 6272: data <= 'd0; 6273: data <= 'd0; 6274: data <= 'd0; 6275: data <= 'd0; 6276: data <= 'd0; 6277: data <= 'd0; 6278: data <= 'd0; 6279: data <= 'd0; 6280: data <= 'd0; 6281: data <= 'd0; 6282: data <= 'd0; 6283: data <= 'd1; 6284: data <= 'd1; 6285: data <= 'd1; 6286: data <= 'd1; 6287: data <= 'd1; 6288: data <= 'd1; 6289: data <= 'd1; 6290: data <= 'd1; 6291: data <= 'd1; 6292: data <= 'd1; 6293: data <= 'd1; 6294: data <= 'd1; 6295: data <= 'd1; 6296: data <= 'd1; 6297: data <= 'd1; 6298: data <= 'd1; 6299: data <= 'd0; 6300: data <= 'd0; 6301: data <= 'd0; 6302: data <= 'd0; 6303: data <= 'd0; 6304: data <= 'd0; 6305: data <= 'd0; 6306: data <= 'd0; 6307: data <= 'd0; 6308: data <= 'd0; 6309: data <= 'd0; 6310: data <= 'd0; 6311: data <= 'd0; 6312: data <= 'd0; 6313: data <= 'd0; 6314: data <= 'd0; 6315: data <= 'd0; 6316: data <= 'd0; 6317: data <= 'd0; 6318: data <= 'd0; 6319: data <= 'd0; 6320: data <= 'd0; 6321: data <= 'd0; 6322: data <= 'd0; 6323: data <= 'd1; 6324: data <= 'd1; 6325: data <= 'd1; 6326: data <= 'd1; 6327: data <= 'd0; 6328: data <= 'd0; 6329: data <= 'd0; 6330: data <= 'd0; 6331: data <= 'd0; 6332: data <= 'd0; 6333: data <= 'd0; 6334: data <= 'd0; 6335: data <= 'd0; 6336: data <= 'd0; 6337: data <= 'd0; 6338: data <= 'd0; 6339: data <= 'd0; 6340: data <= 'd0; 6341: data <= 'd0; 6342: data <= 'd0; 6343: data <= 'd0; 6344: data <= 'd0; 6345: data <= 'd0; 6346: data <= 'd0; 6347: data <= 'd0; 6348: data <= 'd0; 6349: data <= 'd0; 6350: data <= 'd0; 6351: data <= 'd0; 6352: data <= 'd0; 6353: data <= 'd0; 6354: data <= 'd0; 6355: data <= 'd0; 6356: data <= 'd0; 6357: data <= 'd0; 6358: data <= 'd0; 6359: data <= 'd0; 6360: data <= 'd0; 6361: data <= 'd0; 6362: data <= 'd0; 6363: data <= 'd0; 6364: data <= 'd0; 6365: data <= 'd0; 6366: data <= 'd0; 6367: data <= 'd0; 6368: data <= 'd0; 6369: data <= 'd0; 6370: data <= 'd0; 6371: data <= 'd0; 6372: data <= 'd0; 6373: data <= 'd0; 6374: data <= 'd0; 6375: data <= 'd0; 6376: data <= 'd0; 6377: data <= 'd0; 6378: data <= 'd0; 6379: data <= 'd0; 6380: data <= 'd0; 6381: data <= 'd0; 6382: data <= 'd0; 6383: data <= 'd0; 6384: data <= 'd0; 6385: data <= 'd0; 6386: data <= 'd0; 6387: data <= 'd0; 6388: data <= 'd0; 6389: data <= 'd0; 6390: data <= 'd0; 6391: data <= 'd0; 6392: data <= 'd0; 6393: data <= 'd0; 6394: data <= 'd0; 6395: data <= 'd0; 6396: data <= 'd0; 6397: data <= 'd0; 6398: data <= 'd0; 6399: data <= 'd0; 6400: data <= 'd0; 6401: data <= 'd0; 6402: data <= 'd0; 6403: data <= 'd0; 6404: data <= 'd0; 6405: data <= 'd0; 6406: data <= 'd0; 6407: data <= 'd0; 6408: data <= 'd0; 6409: data <= 'd0; 6410: data <= 'd1; 6411: data <= 'd1; 6412: data <= 'd1; 6413: data <= 'd1; 6414: data <= 'd1; 6415: data <= 'd1; 6416: data <= 'd1; 6417: data <= 'd1; 6418: data <= 'd0; 6419: data <= 'd0; 6420: data <= 'd0; 6421: data <= 'd0; 6422: data <= 'd1; 6423: data <= 'd1; 6424: data <= 'd1; 6425: data <= 'd1; 6426: data <= 'd1; 6427: data <= 'd0; 6428: data <= 'd0; 6429: data <= 'd0; 6430: data <= 'd0; 6431: data <= 'd0; 6432: data <= 'd0; 6433: data <= 'd0; 6434: data <= 'd0; 6435: data <= 'd0; 6436: data <= 'd0; 6437: data <= 'd0; 6438: data <= 'd0; 6439: data <= 'd0; 6440: data <= 'd0; 6441: data <= 'd0; 6442: data <= 'd0; 6443: data <= 'd0; 6444: data <= 'd0; 6445: data <= 'd0; 6446: data <= 'd0; 6447: data <= 'd0; 6448: data <= 'd0; 6449: data <= 'd0; 6450: data <= 'd0; 6451: data <= 'd1; 6452: data <= 'd1; 6453: data <= 'd1; 6454: data <= 'd0; 6455: data <= 'd0; 6456: data <= 'd0; 6457: data <= 'd0; 6458: data <= 'd0; 6459: data <= 'd0; 6460: data <= 'd0; 6461: data <= 'd0; 6462: data <= 'd0; 6463: data <= 'd0; 6464: data <= 'd0; 6465: data <= 'd0; 6466: data <= 'd0; 6467: data <= 'd0; 6468: data <= 'd0; 6469: data <= 'd0; 6470: data <= 'd0; 6471: data <= 'd0; 6472: data <= 'd0; 6473: data <= 'd0; 6474: data <= 'd0; 6475: data <= 'd0; 6476: data <= 'd0; 6477: data <= 'd0; 6478: data <= 'd0; 6479: data <= 'd0; 6480: data <= 'd0; 6481: data <= 'd0; 6482: data <= 'd0; 6483: data <= 'd0; 6484: data <= 'd0; 6485: data <= 'd0; 6486: data <= 'd0; 6487: data <= 'd0; 6488: data <= 'd0; 6489: data <= 'd0; 6490: data <= 'd0; 6491: data <= 'd0; 6492: data <= 'd0; 6493: data <= 'd0; 6494: data <= 'd0; 6495: data <= 'd0; 6496: data <= 'd0; 6497: data <= 'd0; 6498: data <= 'd0; 6499: data <= 'd0; 6500: data <= 'd0; 6501: data <= 'd0; 6502: data <= 'd0; 6503: data <= 'd0; 6504: data <= 'd0; 6505: data <= 'd0; 6506: data <= 'd0; 6507: data <= 'd0; 6508: data <= 'd0; 6509: data <= 'd0; 6510: data <= 'd0; 6511: data <= 'd0; 6512: data <= 'd0; 6513: data <= 'd0; 6514: data <= 'd0; 6515: data <= 'd0; 6516: data <= 'd0; 6517: data <= 'd0; 6518: data <= 'd0; 6519: data <= 'd0; 6520: data <= 'd0; 6521: data <= 'd0; 6522: data <= 'd0; 6523: data <= 'd0; 6524: data <= 'd0; 6525: data <= 'd0; 6526: data <= 'd0; 6527: data <= 'd0; 6528: data <= 'd0; 6529: data <= 'd0; 6530: data <= 'd0; 6531: data <= 'd0; 6532: data <= 'd0; 6533: data <= 'd0; 6534: data <= 'd0; 6535: data <= 'd0; 6536: data <= 'd0; 6537: data <= 'd0; 6538: data <= 'd1; 6539: data <= 'd1; 6540: data <= 'd1; 6541: data <= 'd1; 6542: data <= 'd1; 6543: data <= 'd1; 6544: data <= 'd1; 6545: data <= 'd0; 6546: data <= 'd0; 6547: data <= 'd0; 6548: data <= 'd0; 6549: data <= 'd0; 6550: data <= 'd0; 6551: data <= 'd1; 6552: data <= 'd1; 6553: data <= 'd1; 6554: data <= 'd1; 6555: data <= 'd0; 6556: data <= 'd0; 6557: data <= 'd0; 6558: data <= 'd0; 6559: data <= 'd0; 6560: data <= 'd0; 6561: data <= 'd0; 6562: data <= 'd0; 6563: data <= 'd0; 6564: data <= 'd0; 6565: data <= 'd0; 6566: data <= 'd0; 6567: data <= 'd0; 6568: data <= 'd0; 6569: data <= 'd0; 6570: data <= 'd0; 6571: data <= 'd0; 6572: data <= 'd0; 6573: data <= 'd0; 6574: data <= 'd0; 6575: data <= 'd0; 6576: data <= 'd0; 6577: data <= 'd0; 6578: data <= 'd0; 6579: data <= 'd1; 6580: data <= 'd1; 6581: data <= 'd0; 6582: data <= 'd0; 6583: data <= 'd0; 6584: data <= 'd0; 6585: data <= 'd0; 6586: data <= 'd0; 6587: data <= 'd0; 6588: data <= 'd0; 6589: data <= 'd0; 6590: data <= 'd0; 6591: data <= 'd0; 6592: data <= 'd0; 6593: data <= 'd0; 6594: data <= 'd0; 6595: data <= 'd0; 6596: data <= 'd0; 6597: data <= 'd0; 6598: data <= 'd0; 6599: data <= 'd0; 6600: data <= 'd0; 6601: data <= 'd0; 6602: data <= 'd0; 6603: data <= 'd0; 6604: data <= 'd0; 6605: data <= 'd0; 6606: data <= 'd0; 6607: data <= 'd0; 6608: data <= 'd0; 6609: data <= 'd0; 6610: data <= 'd0; 6611: data <= 'd0; 6612: data <= 'd0; 6613: data <= 'd0; 6614: data <= 'd0; 6615: data <= 'd0; 6616: data <= 'd0; 6617: data <= 'd0; 6618: data <= 'd0; 6619: data <= 'd0; 6620: data <= 'd0; 6621: data <= 'd0; 6622: data <= 'd0; 6623: data <= 'd0; 6624: data <= 'd0; 6625: data <= 'd0; 6626: data <= 'd0; 6627: data <= 'd0; 6628: data <= 'd0; 6629: data <= 'd0; 6630: data <= 'd0; 6631: data <= 'd0; 6632: data <= 'd0; 6633: data <= 'd0; 6634: data <= 'd0; 6635: data <= 'd0; 6636: data <= 'd0; 6637: data <= 'd0; 6638: data <= 'd0; 6639: data <= 'd0; 6640: data <= 'd0; 6641: data <= 'd0; 6642: data <= 'd0; 6643: data <= 'd0; 6644: data <= 'd0; 6645: data <= 'd0; 6646: data <= 'd0; 6647: data <= 'd0; 6648: data <= 'd0; 6649: data <= 'd0; 6650: data <= 'd0; 6651: data <= 'd0; 6652: data <= 'd0; 6653: data <= 'd0; 6654: data <= 'd0; 6655: data <= 'd0; 6656: data <= 'd0; 6657: data <= 'd0; 6658: data <= 'd0; 6659: data <= 'd0; 6660: data <= 'd0; 6661: data <= 'd0; 6662: data <= 'd0; 6663: data <= 'd0; 6664: data <= 'd0; 6665: data <= 'd1; 6666: data <= 'd1; 6667: data <= 'd1; 6668: data <= 'd1; 6669: data <= 'd1; 6670: data <= 'd1; 6671: data <= 'd1; 6672: data <= 'd0; 6673: data <= 'd0; 6674: data <= 'd0; 6675: data <= 'd0; 6676: data <= 'd0; 6677: data <= 'd0; 6678: data <= 'd0; 6679: data <= 'd0; 6680: data <= 'd1; 6681: data <= 'd1; 6682: data <= 'd1; 6683: data <= 'd0; 6684: data <= 'd0; 6685: data <= 'd0; 6686: data <= 'd0; 6687: data <= 'd0; 6688: data <= 'd0; 6689: data <= 'd0; 6690: data <= 'd0; 6691: data <= 'd0; 6692: data <= 'd0; 6693: data <= 'd0; 6694: data <= 'd0; 6695: data <= 'd0; 6696: data <= 'd0; 6697: data <= 'd0; 6698: data <= 'd0; 6699: data <= 'd0; 6700: data <= 'd0; 6701: data <= 'd0; 6702: data <= 'd0; 6703: data <= 'd0; 6704: data <= 'd0; 6705: data <= 'd0; 6706: data <= 'd0; 6707: data <= 'd1; 6708: data <= 'd1; 6709: data <= 'd0; 6710: data <= 'd0; 6711: data <= 'd0; 6712: data <= 'd0; 6713: data <= 'd0; 6714: data <= 'd0; 6715: data <= 'd0; 6716: data <= 'd0; 6717: data <= 'd0; 6718: data <= 'd0; 6719: data <= 'd0; 6720: data <= 'd0; 6721: data <= 'd0; 6722: data <= 'd0; 6723: data <= 'd0; 6724: data <= 'd0; 6725: data <= 'd0; 6726: data <= 'd0; 6727: data <= 'd0; 6728: data <= 'd0; 6729: data <= 'd0; 6730: data <= 'd0; 6731: data <= 'd0; 6732: data <= 'd0; 6733: data <= 'd0; 6734: data <= 'd0; 6735: data <= 'd0; 6736: data <= 'd0; 6737: data <= 'd0; 6738: data <= 'd0; 6739: data <= 'd0; 6740: data <= 'd0; 6741: data <= 'd0; 6742: data <= 'd0; 6743: data <= 'd0; 6744: data <= 'd0; 6745: data <= 'd0; 6746: data <= 'd0; 6747: data <= 'd0; 6748: data <= 'd0; 6749: data <= 'd0; 6750: data <= 'd0; 6751: data <= 'd0; 6752: data <= 'd0; 6753: data <= 'd0; 6754: data <= 'd0; 6755: data <= 'd0; 6756: data <= 'd0; 6757: data <= 'd0; 6758: data <= 'd0; 6759: data <= 'd0; 6760: data <= 'd0; 6761: data <= 'd0; 6762: data <= 'd0; 6763: data <= 'd0; 6764: data <= 'd0; 6765: data <= 'd0; 6766: data <= 'd0; 6767: data <= 'd0; 6768: data <= 'd0; 6769: data <= 'd0; 6770: data <= 'd0; 6771: data <= 'd0; 6772: data <= 'd0; 6773: data <= 'd0; 6774: data <= 'd0; 6775: data <= 'd0; 6776: data <= 'd0; 6777: data <= 'd0; 6778: data <= 'd0; 6779: data <= 'd0; 6780: data <= 'd0; 6781: data <= 'd0; 6782: data <= 'd0; 6783: data <= 'd0; 6784: data <= 'd0; 6785: data <= 'd0; 6786: data <= 'd0; 6787: data <= 'd0; 6788: data <= 'd0; 6789: data <= 'd0; 6790: data <= 'd0; 6791: data <= 'd0; 6792: data <= 'd0; 6793: data <= 'd1; 6794: data <= 'd1; 6795: data <= 'd1; 6796: data <= 'd1; 6797: data <= 'd1; 6798: data <= 'd1; 6799: data <= 'd0; 6800: data <= 'd0; 6801: data <= 'd0; 6802: data <= 'd0; 6803: data <= 'd0; 6804: data <= 'd0; 6805: data <= 'd0; 6806: data <= 'd0; 6807: data <= 'd0; 6808: data <= 'd1; 6809: data <= 'd1; 6810: data <= 'd1; 6811: data <= 'd0; 6812: data <= 'd0; 6813: data <= 'd0; 6814: data <= 'd0; 6815: data <= 'd0; 6816: data <= 'd0; 6817: data <= 'd0; 6818: data <= 'd0; 6819: data <= 'd0; 6820: data <= 'd0; 6821: data <= 'd0; 6822: data <= 'd0; 6823: data <= 'd0; 6824: data <= 'd0; 6825: data <= 'd0; 6826: data <= 'd0; 6827: data <= 'd0; 6828: data <= 'd0; 6829: data <= 'd0; 6830: data <= 'd0; 6831: data <= 'd0; 6832: data <= 'd0; 6833: data <= 'd0; 6834: data <= 'd0; 6835: data <= 'd0; 6836: data <= 'd0; 6837: data <= 'd0; 6838: data <= 'd0; 6839: data <= 'd0; 6840: data <= 'd0; 6841: data <= 'd0; 6842: data <= 'd0; 6843: data <= 'd0; 6844: data <= 'd0; 6845: data <= 'd0; 6846: data <= 'd0; 6847: data <= 'd0; 6848: data <= 'd0; 6849: data <= 'd0; 6850: data <= 'd0; 6851: data <= 'd0; 6852: data <= 'd0; 6853: data <= 'd0; 6854: data <= 'd0; 6855: data <= 'd0; 6856: data <= 'd0; 6857: data <= 'd0; 6858: data <= 'd0; 6859: data <= 'd0; 6860: data <= 'd0; 6861: data <= 'd0; 6862: data <= 'd0; 6863: data <= 'd0; 6864: data <= 'd0; 6865: data <= 'd0; 6866: data <= 'd0; 6867: data <= 'd0; 6868: data <= 'd0; 6869: data <= 'd0; 6870: data <= 'd0; 6871: data <= 'd0; 6872: data <= 'd0; 6873: data <= 'd0; 6874: data <= 'd0; 6875: data <= 'd0; 6876: data <= 'd0; 6877: data <= 'd0; 6878: data <= 'd0; 6879: data <= 'd0; 6880: data <= 'd0; 6881: data <= 'd0; 6882: data <= 'd0; 6883: data <= 'd0; 6884: data <= 'd0; 6885: data <= 'd0; 6886: data <= 'd0; 6887: data <= 'd0; 6888: data <= 'd0; 6889: data <= 'd0; 6890: data <= 'd0; 6891: data <= 'd0; 6892: data <= 'd0; 6893: data <= 'd0; 6894: data <= 'd0; 6895: data <= 'd0; 6896: data <= 'd0; 6897: data <= 'd0; 6898: data <= 'd0; 6899: data <= 'd0; 6900: data <= 'd0; 6901: data <= 'd0; 6902: data <= 'd0; 6903: data <= 'd0; 6904: data <= 'd0; 6905: data <= 'd0; 6906: data <= 'd0; 6907: data <= 'd0; 6908: data <= 'd0; 6909: data <= 'd0; 6910: data <= 'd0; 6911: data <= 'd0; 6912: data <= 'd0; 6913: data <= 'd0; 6914: data <= 'd0; 6915: data <= 'd0; 6916: data <= 'd0; 6917: data <= 'd0; 6918: data <= 'd0; 6919: data <= 'd0; 6920: data <= 'd0; 6921: data <= 'd1; 6922: data <= 'd1; 6923: data <= 'd1; 6924: data <= 'd1; 6925: data <= 'd1; 6926: data <= 'd0; 6927: data <= 'd0; 6928: data <= 'd0; 6929: data <= 'd0; 6930: data <= 'd0; 6931: data <= 'd0; 6932: data <= 'd0; 6933: data <= 'd0; 6934: data <= 'd0; 6935: data <= 'd0; 6936: data <= 'd1; 6937: data <= 'd1; 6938: data <= 'd1; 6939: data <= 'd0; 6940: data <= 'd0; 6941: data <= 'd0; 6942: data <= 'd0; 6943: data <= 'd0; 6944: data <= 'd0; 6945: data <= 'd0; 6946: data <= 'd0; 6947: data <= 'd0; 6948: data <= 'd0; 6949: data <= 'd0; 6950: data <= 'd0; 6951: data <= 'd0; 6952: data <= 'd0; 6953: data <= 'd0; 6954: data <= 'd0; 6955: data <= 'd0; 6956: data <= 'd0; 6957: data <= 'd0; 6958: data <= 'd0; 6959: data <= 'd0; 6960: data <= 'd0; 6961: data <= 'd0; 6962: data <= 'd0; 6963: data <= 'd0; 6964: data <= 'd0; 6965: data <= 'd0; 6966: data <= 'd0; 6967: data <= 'd0; 6968: data <= 'd0; 6969: data <= 'd0; 6970: data <= 'd0; 6971: data <= 'd0; 6972: data <= 'd0; 6973: data <= 'd0; 6974: data <= 'd0; 6975: data <= 'd0; 6976: data <= 'd0; 6977: data <= 'd0; 6978: data <= 'd0; 6979: data <= 'd0; 6980: data <= 'd0; 6981: data <= 'd0; 6982: data <= 'd0; 6983: data <= 'd0; 6984: data <= 'd0; 6985: data <= 'd0; 6986: data <= 'd0; 6987: data <= 'd0; 6988: data <= 'd0; 6989: data <= 'd0; 6990: data <= 'd0; 6991: data <= 'd0; 6992: data <= 'd0; 6993: data <= 'd0; 6994: data <= 'd0; 6995: data <= 'd0; 6996: data <= 'd0; 6997: data <= 'd0; 6998: data <= 'd0; 6999: data <= 'd0; 7000: data <= 'd0; 7001: data <= 'd0; 7002: data <= 'd0; 7003: data <= 'd0; 7004: data <= 'd0; 7005: data <= 'd0; 7006: data <= 'd0; 7007: data <= 'd0; 7008: data <= 'd0; 7009: data <= 'd0; 7010: data <= 'd0; 7011: data <= 'd0; 7012: data <= 'd0; 7013: data <= 'd0; 7014: data <= 'd0; 7015: data <= 'd0; 7016: data <= 'd0; 7017: data <= 'd0; 7018: data <= 'd0; 7019: data <= 'd0; 7020: data <= 'd0; 7021: data <= 'd0; 7022: data <= 'd0; 7023: data <= 'd0; 7024: data <= 'd0; 7025: data <= 'd0; 7026: data <= 'd0; 7027: data <= 'd0; 7028: data <= 'd0; 7029: data <= 'd0; 7030: data <= 'd0; 7031: data <= 'd0; 7032: data <= 'd0; 7033: data <= 'd0; 7034: data <= 'd0; 7035: data <= 'd0; 7036: data <= 'd0; 7037: data <= 'd0; 7038: data <= 'd0; 7039: data <= 'd0; 7040: data <= 'd0; 7041: data <= 'd0; 7042: data <= 'd0; 7043: data <= 'd0; 7044: data <= 'd0; 7045: data <= 'd0; 7046: data <= 'd0; 7047: data <= 'd0; 7048: data <= 'd0; 7049: data <= 'd1; 7050: data <= 'd1; 7051: data <= 'd1; 7052: data <= 'd1; 7053: data <= 'd1; 7054: data <= 'd0; 7055: data <= 'd0; 7056: data <= 'd0; 7057: data <= 'd0; 7058: data <= 'd0; 7059: data <= 'd0; 7060: data <= 'd0; 7061: data <= 'd0; 7062: data <= 'd0; 7063: data <= 'd0; 7064: data <= 'd1; 7065: data <= 'd1; 7066: data <= 'd0; 7067: data <= 'd0; 7068: data <= 'd0; 7069: data <= 'd0; 7070: data <= 'd0; 7071: data <= 'd0; 7072: data <= 'd0; 7073: data <= 'd0; 7074: data <= 'd0; 7075: data <= 'd0; 7076: data <= 'd0; 7077: data <= 'd0; 7078: data <= 'd0; 7079: data <= 'd0; 7080: data <= 'd0; 7081: data <= 'd0; 7082: data <= 'd0; 7083: data <= 'd0; 7084: data <= 'd0; 7085: data <= 'd0; 7086: data <= 'd0; 7087: data <= 'd0; 7088: data <= 'd0; 7089: data <= 'd0; 7090: data <= 'd0; 7091: data <= 'd0; 7092: data <= 'd0; 7093: data <= 'd0; 7094: data <= 'd0; 7095: data <= 'd0; 7096: data <= 'd0; 7097: data <= 'd0; 7098: data <= 'd0; 7099: data <= 'd0; 7100: data <= 'd0; 7101: data <= 'd0; 7102: data <= 'd0; 7103: data <= 'd0; 7104: data <= 'd0; 7105: data <= 'd0; 7106: data <= 'd0; 7107: data <= 'd0; 7108: data <= 'd0; 7109: data <= 'd0; 7110: data <= 'd0; 7111: data <= 'd0; 7112: data <= 'd0; 7113: data <= 'd0; 7114: data <= 'd0; 7115: data <= 'd0; 7116: data <= 'd0; 7117: data <= 'd0; 7118: data <= 'd0; 7119: data <= 'd0; 7120: data <= 'd0; 7121: data <= 'd0; 7122: data <= 'd0; 7123: data <= 'd0; 7124: data <= 'd0; 7125: data <= 'd0; 7126: data <= 'd0; 7127: data <= 'd0; 7128: data <= 'd0; 7129: data <= 'd0; 7130: data <= 'd0; 7131: data <= 'd0; 7132: data <= 'd0; 7133: data <= 'd0; 7134: data <= 'd0; 7135: data <= 'd0; 7136: data <= 'd0; 7137: data <= 'd0; 7138: data <= 'd0; 7139: data <= 'd0; 7140: data <= 'd0; 7141: data <= 'd0; 7142: data <= 'd0; 7143: data <= 'd0; 7144: data <= 'd0; 7145: data <= 'd0; 7146: data <= 'd0; 7147: data <= 'd0; 7148: data <= 'd0; 7149: data <= 'd0; 7150: data <= 'd0; 7151: data <= 'd0; 7152: data <= 'd0; 7153: data <= 'd0; 7154: data <= 'd0; 7155: data <= 'd0; 7156: data <= 'd0; 7157: data <= 'd0; 7158: data <= 'd0; 7159: data <= 'd0; 7160: data <= 'd0; 7161: data <= 'd0; 7162: data <= 'd0; 7163: data <= 'd0; 7164: data <= 'd0; 7165: data <= 'd0; 7166: data <= 'd0; 7167: data <= 'd0; 7168: data <= 'd0; 7169: data <= 'd0; 7170: data <= 'd0; 7171: data <= 'd0; 7172: data <= 'd0; 7173: data <= 'd0; 7174: data <= 'd0; 7175: data <= 'd0; 7176: data <= 'd1; 7177: data <= 'd1; 7178: data <= 'd1; 7179: data <= 'd1; 7180: data <= 'd1; 7181: data <= 'd1; 7182: data <= 'd0; 7183: data <= 'd0; 7184: data <= 'd0; 7185: data <= 'd0; 7186: data <= 'd0; 7187: data <= 'd0; 7188: data <= 'd0; 7189: data <= 'd0; 7190: data <= 'd0; 7191: data <= 'd0; 7192: data <= 'd0; 7193: data <= 'd0; 7194: data <= 'd0; 7195: data <= 'd0; 7196: data <= 'd0; 7197: data <= 'd0; 7198: data <= 'd0; 7199: data <= 'd0; 7200: data <= 'd0; 7201: data <= 'd0; 7202: data <= 'd0; 7203: data <= 'd0; 7204: data <= 'd0; 7205: data <= 'd0; 7206: data <= 'd0; 7207: data <= 'd0; 7208: data <= 'd0; 7209: data <= 'd0; 7210: data <= 'd0; 7211: data <= 'd0; 7212: data <= 'd0; 7213: data <= 'd0; 7214: data <= 'd0; 7215: data <= 'd0; 7216: data <= 'd0; 7217: data <= 'd0; 7218: data <= 'd0; 7219: data <= 'd0; 7220: data <= 'd0; 7221: data <= 'd0; 7222: data <= 'd0; 7223: data <= 'd0; 7224: data <= 'd0; 7225: data <= 'd0; 7226: data <= 'd0; 7227: data <= 'd0; 7228: data <= 'd0; 7229: data <= 'd0; 7230: data <= 'd0; 7231: data <= 'd0; 7232: data <= 'd0; 7233: data <= 'd0; 7234: data <= 'd0; 7235: data <= 'd0; 7236: data <= 'd0; 7237: data <= 'd0; 7238: data <= 'd0; 7239: data <= 'd0; 7240: data <= 'd0; 7241: data <= 'd0; 7242: data <= 'd0; 7243: data <= 'd0; 7244: data <= 'd0; 7245: data <= 'd0; 7246: data <= 'd0; 7247: data <= 'd0; 7248: data <= 'd0; 7249: data <= 'd0; 7250: data <= 'd0; 7251: data <= 'd0; 7252: data <= 'd0; 7253: data <= 'd0; 7254: data <= 'd0; 7255: data <= 'd0; 7256: data <= 'd0; 7257: data <= 'd0; 7258: data <= 'd0; 7259: data <= 'd0; 7260: data <= 'd0; 7261: data <= 'd0; 7262: data <= 'd0; 7263: data <= 'd0; 7264: data <= 'd0; 7265: data <= 'd0; 7266: data <= 'd0; 7267: data <= 'd0; 7268: data <= 'd0; 7269: data <= 'd0; 7270: data <= 'd0; 7271: data <= 'd0; 7272: data <= 'd0; 7273: data <= 'd0; 7274: data <= 'd0; 7275: data <= 'd0; 7276: data <= 'd0; 7277: data <= 'd0; 7278: data <= 'd0; 7279: data <= 'd0; 7280: data <= 'd0; 7281: data <= 'd0; 7282: data <= 'd0; 7283: data <= 'd0; 7284: data <= 'd0; 7285: data <= 'd0; 7286: data <= 'd0; 7287: data <= 'd0; 7288: data <= 'd0; 7289: data <= 'd0; 7290: data <= 'd0; 7291: data <= 'd0; 7292: data <= 'd0; 7293: data <= 'd0; 7294: data <= 'd0; 7295: data <= 'd0; 7296: data <= 'd0; 7297: data <= 'd0; 7298: data <= 'd0; 7299: data <= 'd0; 7300: data <= 'd0; 7301: data <= 'd0; 7302: data <= 'd0; 7303: data <= 'd0; 7304: data <= 'd1; 7305: data <= 'd1; 7306: data <= 'd1; 7307: data <= 'd1; 7308: data <= 'd1; 7309: data <= 'd0; 7310: data <= 'd0; 7311: data <= 'd0; 7312: data <= 'd0; 7313: data <= 'd0; 7314: data <= 'd0; 7315: data <= 'd0; 7316: data <= 'd0; 7317: data <= 'd0; 7318: data <= 'd0; 7319: data <= 'd0; 7320: data <= 'd0; 7321: data <= 'd0; 7322: data <= 'd0; 7323: data <= 'd0; 7324: data <= 'd0; 7325: data <= 'd0; 7326: data <= 'd0; 7327: data <= 'd0; 7328: data <= 'd0; 7329: data <= 'd0; 7330: data <= 'd0; 7331: data <= 'd0; 7332: data <= 'd0; 7333: data <= 'd0; 7334: data <= 'd0; 7335: data <= 'd0; 7336: data <= 'd0; 7337: data <= 'd0; 7338: data <= 'd0; 7339: data <= 'd0; 7340: data <= 'd0; 7341: data <= 'd0; 7342: data <= 'd0; 7343: data <= 'd0; 7344: data <= 'd0; 7345: data <= 'd0; 7346: data <= 'd0; 7347: data <= 'd0; 7348: data <= 'd0; 7349: data <= 'd0; 7350: data <= 'd0; 7351: data <= 'd0; 7352: data <= 'd0; 7353: data <= 'd0; 7354: data <= 'd0; 7355: data <= 'd0; 7356: data <= 'd0; 7357: data <= 'd0; 7358: data <= 'd0; 7359: data <= 'd0; 7360: data <= 'd0; 7361: data <= 'd0; 7362: data <= 'd0; 7363: data <= 'd0; 7364: data <= 'd0; 7365: data <= 'd0; 7366: data <= 'd0; 7367: data <= 'd0; 7368: data <= 'd0; 7369: data <= 'd0; 7370: data <= 'd0; 7371: data <= 'd0; 7372: data <= 'd0; 7373: data <= 'd0; 7374: data <= 'd0; 7375: data <= 'd0; 7376: data <= 'd0; 7377: data <= 'd0; 7378: data <= 'd0; 7379: data <= 'd0; 7380: data <= 'd0; 7381: data <= 'd0; 7382: data <= 'd0; 7383: data <= 'd0; 7384: data <= 'd0; 7385: data <= 'd0; 7386: data <= 'd0; 7387: data <= 'd0; 7388: data <= 'd0; 7389: data <= 'd0; 7390: data <= 'd0; 7391: data <= 'd0; 7392: data <= 'd0; 7393: data <= 'd0; 7394: data <= 'd0; 7395: data <= 'd0; 7396: data <= 'd0; 7397: data <= 'd0; 7398: data <= 'd0; 7399: data <= 'd0; 7400: data <= 'd0; 7401: data <= 'd0; 7402: data <= 'd0; 7403: data <= 'd0; 7404: data <= 'd0; 7405: data <= 'd0; 7406: data <= 'd0; 7407: data <= 'd0; 7408: data <= 'd0; 7409: data <= 'd0; 7410: data <= 'd0; 7411: data <= 'd0; 7412: data <= 'd0; 7413: data <= 'd0; 7414: data <= 'd0; 7415: data <= 'd0; 7416: data <= 'd0; 7417: data <= 'd0; 7418: data <= 'd0; 7419: data <= 'd0; 7420: data <= 'd0; 7421: data <= 'd0; 7422: data <= 'd0; 7423: data <= 'd0; 7424: data <= 'd0; 7425: data <= 'd0; 7426: data <= 'd0; 7427: data <= 'd0; 7428: data <= 'd0; 7429: data <= 'd0; 7430: data <= 'd0; 7431: data <= 'd1; 7432: data <= 'd1; 7433: data <= 'd1; 7434: data <= 'd1; 7435: data <= 'd1; 7436: data <= 'd1; 7437: data <= 'd0; 7438: data <= 'd0; 7439: data <= 'd0; 7440: data <= 'd0; 7441: data <= 'd0; 7442: data <= 'd0; 7443: data <= 'd0; 7444: data <= 'd0; 7445: data <= 'd0; 7446: data <= 'd0; 7447: data <= 'd0; 7448: data <= 'd0; 7449: data <= 'd0; 7450: data <= 'd0; 7451: data <= 'd0; 7452: data <= 'd0; 7453: data <= 'd0; 7454: data <= 'd0; 7455: data <= 'd0; 7456: data <= 'd0; 7457: data <= 'd0; 7458: data <= 'd0; 7459: data <= 'd0; 7460: data <= 'd0; 7461: data <= 'd0; 7462: data <= 'd0; 7463: data <= 'd0; 7464: data <= 'd0; 7465: data <= 'd0; 7466: data <= 'd0; 7467: data <= 'd0; 7468: data <= 'd0; 7469: data <= 'd0; 7470: data <= 'd0; 7471: data <= 'd0; 7472: data <= 'd0; 7473: data <= 'd0; 7474: data <= 'd0; 7475: data <= 'd0; 7476: data <= 'd0; 7477: data <= 'd0; 7478: data <= 'd0; 7479: data <= 'd0; 7480: data <= 'd0; 7481: data <= 'd0; 7482: data <= 'd0; 7483: data <= 'd0; 7484: data <= 'd0; 7485: data <= 'd0; 7486: data <= 'd0; 7487: data <= 'd0; 7488: data <= 'd0; 7489: data <= 'd0; 7490: data <= 'd0; 7491: data <= 'd0; 7492: data <= 'd0; 7493: data <= 'd0; 7494: data <= 'd0; 7495: data <= 'd0; 7496: data <= 'd0; 7497: data <= 'd0; 7498: data <= 'd0; 7499: data <= 'd0; 7500: data <= 'd0; 7501: data <= 'd0; 7502: data <= 'd0; 7503: data <= 'd0; 7504: data <= 'd0; 7505: data <= 'd0; 7506: data <= 'd0; 7507: data <= 'd0; 7508: data <= 'd0; 7509: data <= 'd0; 7510: data <= 'd0; 7511: data <= 'd0; 7512: data <= 'd0; 7513: data <= 'd0; 7514: data <= 'd0; 7515: data <= 'd0; 7516: data <= 'd0; 7517: data <= 'd0; 7518: data <= 'd0; 7519: data <= 'd0; 7520: data <= 'd0; 7521: data <= 'd0; 7522: data <= 'd0; 7523: data <= 'd0; 7524: data <= 'd0; 7525: data <= 'd0; 7526: data <= 'd0; 7527: data <= 'd0; 7528: data <= 'd0; 7529: data <= 'd0; 7530: data <= 'd0; 7531: data <= 'd0; 7532: data <= 'd0; 7533: data <= 'd0; 7534: data <= 'd0; 7535: data <= 'd0; 7536: data <= 'd0; 7537: data <= 'd0; 7538: data <= 'd0; 7539: data <= 'd0; 7540: data <= 'd0; 7541: data <= 'd0; 7542: data <= 'd0; 7543: data <= 'd0; 7544: data <= 'd0; 7545: data <= 'd0; 7546: data <= 'd0; 7547: data <= 'd0; 7548: data <= 'd0; 7549: data <= 'd0; 7550: data <= 'd0; 7551: data <= 'd0; 7552: data <= 'd0; 7553: data <= 'd1; 7554: data <= 'd1; 7555: data <= 'd0; 7556: data <= 'd0; 7557: data <= 'd0; 7558: data <= 'd0; 7559: data <= 'd1; 7560: data <= 'd1; 7561: data <= 'd1; 7562: data <= 'd1; 7563: data <= 'd1; 7564: data <= 'd1; 7565: data <= 'd1; 7566: data <= 'd0; 7567: data <= 'd0; 7568: data <= 'd0; 7569: data <= 'd0; 7570: data <= 'd0; 7571: data <= 'd0; 7572: data <= 'd0; 7573: data <= 'd0; 7574: data <= 'd0; 7575: data <= 'd0; 7576: data <= 'd0; 7577: data <= 'd0; 7578: data <= 'd0; 7579: data <= 'd0; 7580: data <= 'd0; 7581: data <= 'd0; 7582: data <= 'd0; 7583: data <= 'd0; 7584: data <= 'd0; 7585: data <= 'd0; 7586: data <= 'd0; 7587: data <= 'd0; 7588: data <= 'd0; 7589: data <= 'd0; 7590: data <= 'd0; 7591: data <= 'd0; 7592: data <= 'd0; 7593: data <= 'd0; 7594: data <= 'd0; 7595: data <= 'd0; 7596: data <= 'd0; 7597: data <= 'd0; 7598: data <= 'd0; 7599: data <= 'd0; 7600: data <= 'd0; 7601: data <= 'd0; 7602: data <= 'd0; 7603: data <= 'd0; 7604: data <= 'd0; 7605: data <= 'd0; 7606: data <= 'd0; 7607: data <= 'd0; 7608: data <= 'd0; 7609: data <= 'd0; 7610: data <= 'd0; 7611: data <= 'd0; 7612: data <= 'd0; 7613: data <= 'd0; 7614: data <= 'd0; 7615: data <= 'd0; 7616: data <= 'd0; 7617: data <= 'd0; 7618: data <= 'd0; 7619: data <= 'd0; 7620: data <= 'd0; 7621: data <= 'd0; 7622: data <= 'd0; 7623: data <= 'd0; 7624: data <= 'd0; 7625: data <= 'd0; 7626: data <= 'd0; 7627: data <= 'd0; 7628: data <= 'd0; 7629: data <= 'd0; 7630: data <= 'd0; 7631: data <= 'd0; 7632: data <= 'd0; 7633: data <= 'd0; 7634: data <= 'd0; 7635: data <= 'd0; 7636: data <= 'd0; 7637: data <= 'd0; 7638: data <= 'd0; 7639: data <= 'd0; 7640: data <= 'd0; 7641: data <= 'd0; 7642: data <= 'd0; 7643: data <= 'd0; 7644: data <= 'd0; 7645: data <= 'd0; 7646: data <= 'd0; 7647: data <= 'd0; 7648: data <= 'd0; 7649: data <= 'd0; 7650: data <= 'd0; 7651: data <= 'd0; 7652: data <= 'd0; 7653: data <= 'd0; 7654: data <= 'd0; 7655: data <= 'd0; 7656: data <= 'd0; 7657: data <= 'd0; 7658: data <= 'd0; 7659: data <= 'd0; 7660: data <= 'd0; 7661: data <= 'd0; 7662: data <= 'd0; 7663: data <= 'd0; 7664: data <= 'd0; 7665: data <= 'd0; 7666: data <= 'd0; 7667: data <= 'd0; 7668: data <= 'd0; 7669: data <= 'd0; 7670: data <= 'd0; 7671: data <= 'd0; 7672: data <= 'd0; 7673: data <= 'd0; 7674: data <= 'd0; 7675: data <= 'd0; 7676: data <= 'd0; 7677: data <= 'd0; 7678: data <= 'd0; 7679: data <= 'd0; 7680: data <= 'd0; 7681: data <= 'd0; 7682: data <= 'd1; 7683: data <= 'd1; 7684: data <= 'd0; 7685: data <= 'd1; 7686: data <= 'd1; 7687: data <= 'd1; 7688: data <= 'd1; 7689: data <= 'd1; 7690: data <= 'd1; 7691: data <= 'd1; 7692: data <= 'd1; 7693: data <= 'd1; 7694: data <= 'd0; 7695: data <= 'd0; 7696: data <= 'd0; 7697: data <= 'd0; 7698: data <= 'd0; 7699: data <= 'd0; 7700: data <= 'd0; 7701: data <= 'd0; 7702: data <= 'd0; 7703: data <= 'd0; 7704: data <= 'd0; 7705: data <= 'd0; 7706: data <= 'd0; 7707: data <= 'd0; 7708: data <= 'd0; 7709: data <= 'd0; 7710: data <= 'd0; 7711: data <= 'd0; 7712: data <= 'd0; 7713: data <= 'd0; 7714: data <= 'd0; 7715: data <= 'd0; 7716: data <= 'd0; 7717: data <= 'd0; 7718: data <= 'd0; 7719: data <= 'd0; 7720: data <= 'd0; 7721: data <= 'd0; 7722: data <= 'd0; 7723: data <= 'd0; 7724: data <= 'd0; 7725: data <= 'd0; 7726: data <= 'd0; 7727: data <= 'd0; 7728: data <= 'd0; 7729: data <= 'd0; 7730: data <= 'd0; 7731: data <= 'd0; 7732: data <= 'd0; 7733: data <= 'd0; 7734: data <= 'd0; 7735: data <= 'd0; 7736: data <= 'd0; 7737: data <= 'd0; 7738: data <= 'd0; 7739: data <= 'd0; 7740: data <= 'd0; 7741: data <= 'd0; 7742: data <= 'd0; 7743: data <= 'd0; 7744: data <= 'd0; 7745: data <= 'd0; 7746: data <= 'd0; 7747: data <= 'd0; 7748: data <= 'd0; 7749: data <= 'd0; 7750: data <= 'd0; 7751: data <= 'd0; 7752: data <= 'd0; 7753: data <= 'd0; 7754: data <= 'd0; 7755: data <= 'd0; 7756: data <= 'd0; 7757: data <= 'd0; 7758: data <= 'd0; 7759: data <= 'd0; 7760: data <= 'd0; 7761: data <= 'd0; 7762: data <= 'd0; 7763: data <= 'd0; 7764: data <= 'd0; 7765: data <= 'd0; 7766: data <= 'd0; 7767: data <= 'd0; 7768: data <= 'd0; 7769: data <= 'd0; 7770: data <= 'd0; 7771: data <= 'd0; 7772: data <= 'd0; 7773: data <= 'd0; 7774: data <= 'd0; 7775: data <= 'd0; 7776: data <= 'd0; 7777: data <= 'd0; 7778: data <= 'd0; 7779: data <= 'd0; 7780: data <= 'd0; 7781: data <= 'd0; 7782: data <= 'd0; 7783: data <= 'd0; 7784: data <= 'd0; 7785: data <= 'd0; 7786: data <= 'd0; 7787: data <= 'd0; 7788: data <= 'd0; 7789: data <= 'd0; 7790: data <= 'd0; 7791: data <= 'd0; 7792: data <= 'd0; 7793: data <= 'd0; 7794: data <= 'd0; 7795: data <= 'd0; 7796: data <= 'd0; 7797: data <= 'd0; 7798: data <= 'd0; 7799: data <= 'd0; 7800: data <= 'd0; 7801: data <= 'd0; 7802: data <= 'd0; 7803: data <= 'd0; 7804: data <= 'd0; 7805: data <= 'd0; 7806: data <= 'd0; 7807: data <= 'd0; 7808: data <= 'd0; 7809: data <= 'd0; 7810: data <= 'd0; 7811: data <= 'd1; 7812: data <= 'd1; 7813: data <= 'd1; 7814: data <= 'd1; 7815: data <= 'd1; 7816: data <= 'd1; 7817: data <= 'd1; 7818: data <= 'd1; 7819: data <= 'd1; 7820: data <= 'd1; 7821: data <= 'd1; 7822: data <= 'd0; 7823: data <= 'd0; 7824: data <= 'd0; 7825: data <= 'd0; 7826: data <= 'd0; 7827: data <= 'd0; 7828: data <= 'd0; 7829: data <= 'd0; 7830: data <= 'd0; 7831: data <= 'd0; 7832: data <= 'd0; 7833: data <= 'd0; 7834: data <= 'd0; 7835: data <= 'd0; 7836: data <= 'd0; 7837: data <= 'd0; 7838: data <= 'd0; 7839: data <= 'd0; 7840: data <= 'd0; 7841: data <= 'd0; 7842: data <= 'd0; 7843: data <= 'd0; 7844: data <= 'd0; 7845: data <= 'd0; 7846: data <= 'd0; 7847: data <= 'd0; 7848: data <= 'd0; 7849: data <= 'd0; 7850: data <= 'd0; 7851: data <= 'd0; 7852: data <= 'd0; 7853: data <= 'd0; 7854: data <= 'd0; 7855: data <= 'd0; 7856: data <= 'd0; 7857: data <= 'd0; 7858: data <= 'd0; 7859: data <= 'd0; 7860: data <= 'd0; 7861: data <= 'd0; 7862: data <= 'd0; 7863: data <= 'd0; 7864: data <= 'd0; 7865: data <= 'd0; 7866: data <= 'd0; 7867: data <= 'd0; 7868: data <= 'd0; 7869: data <= 'd0; 7870: data <= 'd0; 7871: data <= 'd0; 7872: data <= 'd0; 7873: data <= 'd0; 7874: data <= 'd0; 7875: data <= 'd0; 7876: data <= 'd0; 7877: data <= 'd0; 7878: data <= 'd0; 7879: data <= 'd0; 7880: data <= 'd0; 7881: data <= 'd0; 7882: data <= 'd0; 7883: data <= 'd0; 7884: data <= 'd0; 7885: data <= 'd0; 7886: data <= 'd0; 7887: data <= 'd0; 7888: data <= 'd0; 7889: data <= 'd0; 7890: data <= 'd0; 7891: data <= 'd0; 7892: data <= 'd0; 7893: data <= 'd0; 7894: data <= 'd0; 7895: data <= 'd0; 7896: data <= 'd0; 7897: data <= 'd0; 7898: data <= 'd0; 7899: data <= 'd0; 7900: data <= 'd0; 7901: data <= 'd0; 7902: data <= 'd0; 7903: data <= 'd0; 7904: data <= 'd0; 7905: data <= 'd0; 7906: data <= 'd0; 7907: data <= 'd0; 7908: data <= 'd0; 7909: data <= 'd0; 7910: data <= 'd0; 7911: data <= 'd0; 7912: data <= 'd0; 7913: data <= 'd0; 7914: data <= 'd0; 7915: data <= 'd0; 7916: data <= 'd0; 7917: data <= 'd0; 7918: data <= 'd0; 7919: data <= 'd0; 7920: data <= 'd0; 7921: data <= 'd0; 7922: data <= 'd0; 7923: data <= 'd0; 7924: data <= 'd0; 7925: data <= 'd0; 7926: data <= 'd0; 7927: data <= 'd0; 7928: data <= 'd0; 7929: data <= 'd0; 7930: data <= 'd0; 7931: data <= 'd0; 7932: data <= 'd0; 7933: data <= 'd0; 7934: data <= 'd0; 7935: data <= 'd0; 7936: data <= 'd0; 7937: data <= 'd0; 7938: data <= 'd0; 7939: data <= 'd0; 7940: data <= 'd1; 7941: data <= 'd1; 7942: data <= 'd1; 7943: data <= 'd1; 7944: data <= 'd0; 7945: data <= 'd1; 7946: data <= 'd1; 7947: data <= 'd1; 7948: data <= 'd1; 7949: data <= 'd1; 7950: data <= 'd0; 7951: data <= 'd0; 7952: data <= 'd0; 7953: data <= 'd0; 7954: data <= 'd0; 7955: data <= 'd0; 7956: data <= 'd0; 7957: data <= 'd0; 7958: data <= 'd0; 7959: data <= 'd0; 7960: data <= 'd0; 7961: data <= 'd0; 7962: data <= 'd0; 7963: data <= 'd0; 7964: data <= 'd0; 7965: data <= 'd0; 7966: data <= 'd0; 7967: data <= 'd0; 7968: data <= 'd0; 7969: data <= 'd0; 7970: data <= 'd0; 7971: data <= 'd0; 7972: data <= 'd0; 7973: data <= 'd0; 7974: data <= 'd0; 7975: data <= 'd0; 7976: data <= 'd0; 7977: data <= 'd0; 7978: data <= 'd0; 7979: data <= 'd0; 7980: data <= 'd0; 7981: data <= 'd0; 7982: data <= 'd0; 7983: data <= 'd0; 7984: data <= 'd0; 7985: data <= 'd0; 7986: data <= 'd0; 7987: data <= 'd0; 7988: data <= 'd0; 7989: data <= 'd0; 7990: data <= 'd0; 7991: data <= 'd0; 7992: data <= 'd0; 7993: data <= 'd0; 7994: data <= 'd0; 7995: data <= 'd0; 7996: data <= 'd0; 7997: data <= 'd0; 7998: data <= 'd0; 7999: data <= 'd0; 8000: data <= 'd0; 8001: data <= 'd0; 8002: data <= 'd0; 8003: data <= 'd0; 8004: data <= 'd0; 8005: data <= 'd0; 8006: data <= 'd0; 8007: data <= 'd0; 8008: data <= 'd0; 8009: data <= 'd0; 8010: data <= 'd0; 8011: data <= 'd0; 8012: data <= 'd0; 8013: data <= 'd0; 8014: data <= 'd0; 8015: data <= 'd0; 8016: data <= 'd0; 8017: data <= 'd0; 8018: data <= 'd0; 8019: data <= 'd0; 8020: data <= 'd0; 8021: data <= 'd0; 8022: data <= 'd0; 8023: data <= 'd0; 8024: data <= 'd0; 8025: data <= 'd0; 8026: data <= 'd0; 8027: data <= 'd0; 8028: data <= 'd0; 8029: data <= 'd0; 8030: data <= 'd0; 8031: data <= 'd0; 8032: data <= 'd0; 8033: data <= 'd0; 8034: data <= 'd0; 8035: data <= 'd0; 8036: data <= 'd0; 8037: data <= 'd0; 8038: data <= 'd0; 8039: data <= 'd0; 8040: data <= 'd0; 8041: data <= 'd0; 8042: data <= 'd0; 8043: data <= 'd0; 8044: data <= 'd0; 8045: data <= 'd0; 8046: data <= 'd0; 8047: data <= 'd0; 8048: data <= 'd0; 8049: data <= 'd0; 8050: data <= 'd0; 8051: data <= 'd0; 8052: data <= 'd0; 8053: data <= 'd0; 8054: data <= 'd0; 8055: data <= 'd0; 8056: data <= 'd0; 8057: data <= 'd0; 8058: data <= 'd0; 8059: data <= 'd0; 8060: data <= 'd0; 8061: data <= 'd0; 8062: data <= 'd0; 8063: data <= 'd0; 8064: data <= 'd0; 8065: data <= 'd0; 8066: data <= 'd0; 8067: data <= 'd0; 8068: data <= 'd1; 8069: data <= 'd0; 8070: data <= 'd0; 8071: data <= 'd0; 8072: data <= 'd0; 8073: data <= 'd0; 8074: data <= 'd1; 8075: data <= 'd1; 8076: data <= 'd1; 8077: data <= 'd1; 8078: data <= 'd0; 8079: data <= 'd0; 8080: data <= 'd0; 8081: data <= 'd0; 8082: data <= 'd0; 8083: data <= 'd0; 8084: data <= 'd0; 8085: data <= 'd0; 8086: data <= 'd0; 8087: data <= 'd0; 8088: data <= 'd0; 8089: data <= 'd0; 8090: data <= 'd0; 8091: data <= 'd0; 8092: data <= 'd0; 8093: data <= 'd0; 8094: data <= 'd0; 8095: data <= 'd0; 8096: data <= 'd0; 8097: data <= 'd0; 8098: data <= 'd0; 8099: data <= 'd0; 8100: data <= 'd0; 8101: data <= 'd0; 8102: data <= 'd0; 8103: data <= 'd0; 8104: data <= 'd0; 8105: data <= 'd0; 8106: data <= 'd0; 8107: data <= 'd0; 8108: data <= 'd0; 8109: data <= 'd0; 8110: data <= 'd0; 8111: data <= 'd0; 8112: data <= 'd0; 8113: data <= 'd0; 8114: data <= 'd0; 8115: data <= 'd0; 8116: data <= 'd0; 8117: data <= 'd0; 8118: data <= 'd0; 8119: data <= 'd0; 8120: data <= 'd0; 8121: data <= 'd0; 8122: data <= 'd0; 8123: data <= 'd0; 8124: data <= 'd0; 8125: data <= 'd0; 8126: data <= 'd0; 8127: data <= 'd0; 8128: data <= 'd0; 8129: data <= 'd0; 8130: data <= 'd0; 8131: data <= 'd0; 8132: data <= 'd0; 8133: data <= 'd0; 8134: data <= 'd0; 8135: data <= 'd0; 8136: data <= 'd0; 8137: data <= 'd0; 8138: data <= 'd0; 8139: data <= 'd0; 8140: data <= 'd0; 8141: data <= 'd0; 8142: data <= 'd0; 8143: data <= 'd0; 8144: data <= 'd0; 8145: data <= 'd0; 8146: data <= 'd0; 8147: data <= 'd0; 8148: data <= 'd0; 8149: data <= 'd0; 8150: data <= 'd0; 8151: data <= 'd0; 8152: data <= 'd0; 8153: data <= 'd0; 8154: data <= 'd0; 8155: data <= 'd0; 8156: data <= 'd0; 8157: data <= 'd0; 8158: data <= 'd0; 8159: data <= 'd0; 8160: data <= 'd0; 8161: data <= 'd0; 8162: data <= 'd0; 8163: data <= 'd0; 8164: data <= 'd0; 8165: data <= 'd0; 8166: data <= 'd0; 8167: data <= 'd0; 8168: data <= 'd0; 8169: data <= 'd0; 8170: data <= 'd0; 8171: data <= 'd0; 8172: data <= 'd0; 8173: data <= 'd0; 8174: data <= 'd0; 8175: data <= 'd0; 8176: data <= 'd0; 8177: data <= 'd0; 8178: data <= 'd0; 8179: data <= 'd0; 8180: data <= 'd0; 8181: data <= 'd0; 8182: data <= 'd0; 8183: data <= 'd0; 8184: data <= 'd0; 8185: data <= 'd0; 8186: data <= 'd0; 8187: data <= 'd0; 8188: data <= 'd0; 8189: data <= 'd0; 8190: data <= 'd0; 8191: data <= 'd0; 8192: data <= 'd0; 8193: data <= 'd0; 8194: data <= 'd0; 8195: data <= 'd0; 8196: data <= 'd0; 8197: data <= 'd0; 8198: data <= 'd0; 8199: data <= 'd0; 8200: data <= 'd0; 8201: data <= 'd0; 8202: data <= 'd1; 8203: data <= 'd1; 8204: data <= 'd1; 8205: data <= 'd1; 8206: data <= 'd1; 8207: data <= 'd0; 8208: data <= 'd0; 8209: data <= 'd0; 8210: data <= 'd0; 8211: data <= 'd0; 8212: data <= 'd0; 8213: data <= 'd0; 8214: data <= 'd0; 8215: data <= 'd0; 8216: data <= 'd0; 8217: data <= 'd0; 8218: data <= 'd0; 8219: data <= 'd0; 8220: data <= 'd0; 8221: data <= 'd0; 8222: data <= 'd0; 8223: data <= 'd0; 8224: data <= 'd0; 8225: data <= 'd0; 8226: data <= 'd0; 8227: data <= 'd0; 8228: data <= 'd0; 8229: data <= 'd0; 8230: data <= 'd0; 8231: data <= 'd0; 8232: data <= 'd0; 8233: data <= 'd0; 8234: data <= 'd0; 8235: data <= 'd0; 8236: data <= 'd0; 8237: data <= 'd0; 8238: data <= 'd0; 8239: data <= 'd0; 8240: data <= 'd0; 8241: data <= 'd0; 8242: data <= 'd0; 8243: data <= 'd0; 8244: data <= 'd0; 8245: data <= 'd0; 8246: data <= 'd0; 8247: data <= 'd0; 8248: data <= 'd0; 8249: data <= 'd0; 8250: data <= 'd0; 8251: data <= 'd0; 8252: data <= 'd0; 8253: data <= 'd0; 8254: data <= 'd0; 8255: data <= 'd0; 8256: data <= 'd0; 8257: data <= 'd0; 8258: data <= 'd0; 8259: data <= 'd0; 8260: data <= 'd0; 8261: data <= 'd0; 8262: data <= 'd0; 8263: data <= 'd0; 8264: data <= 'd0; 8265: data <= 'd0; 8266: data <= 'd0; 8267: data <= 'd0; 8268: data <= 'd0; 8269: data <= 'd0; 8270: data <= 'd0; 8271: data <= 'd0; 8272: data <= 'd0; 8273: data <= 'd0; 8274: data <= 'd0; 8275: data <= 'd0; 8276: data <= 'd0; 8277: data <= 'd0; 8278: data <= 'd0; 8279: data <= 'd0; 8280: data <= 'd0; 8281: data <= 'd0; 8282: data <= 'd0; 8283: data <= 'd0; 8284: data <= 'd0; 8285: data <= 'd0; 8286: data <= 'd0; 8287: data <= 'd0; 8288: data <= 'd0; 8289: data <= 'd0; 8290: data <= 'd0; 8291: data <= 'd0; 8292: data <= 'd0; 8293: data <= 'd0; 8294: data <= 'd0; 8295: data <= 'd0; 8296: data <= 'd0; 8297: data <= 'd0; 8298: data <= 'd0; 8299: data <= 'd0; 8300: data <= 'd0; 8301: data <= 'd0; 8302: data <= 'd0; 8303: data <= 'd0; 8304: data <= 'd0; 8305: data <= 'd0; 8306: data <= 'd0; 8307: data <= 'd0; 8308: data <= 'd0; 8309: data <= 'd0; 8310: data <= 'd0; 8311: data <= 'd0; 8312: data <= 'd0; 8313: data <= 'd0; 8314: data <= 'd0; 8315: data <= 'd0; 8316: data <= 'd0; 8317: data <= 'd0; 8318: data <= 'd0; 8319: data <= 'd0; 8320: data <= 'd0; 8321: data <= 'd0; 8322: data <= 'd0; 8323: data <= 'd0; 8324: data <= 'd0; 8325: data <= 'd0; 8326: data <= 'd0; 8327: data <= 'd0; 8328: data <= 'd0; 8329: data <= 'd0; 8330: data <= 'd1; 8331: data <= 'd1; 8332: data <= 'd1; 8333: data <= 'd1; 8334: data <= 'd1; 8335: data <= 'd0; 8336: data <= 'd0; 8337: data <= 'd0; 8338: data <= 'd0; 8339: data <= 'd0; 8340: data <= 'd0; 8341: data <= 'd0; 8342: data <= 'd0; 8343: data <= 'd0; 8344: data <= 'd0; 8345: data <= 'd0; 8346: data <= 'd0; 8347: data <= 'd0; 8348: data <= 'd0; 8349: data <= 'd0; 8350: data <= 'd0; 8351: data <= 'd0; 8352: data <= 'd0; 8353: data <= 'd0; 8354: data <= 'd0; 8355: data <= 'd0; 8356: data <= 'd0; 8357: data <= 'd0; 8358: data <= 'd0; 8359: data <= 'd0; 8360: data <= 'd0; 8361: data <= 'd0; 8362: data <= 'd0; 8363: data <= 'd0; 8364: data <= 'd0; 8365: data <= 'd0; 8366: data <= 'd0; 8367: data <= 'd0; 8368: data <= 'd0; 8369: data <= 'd0; 8370: data <= 'd0; 8371: data <= 'd0; 8372: data <= 'd0; 8373: data <= 'd0; 8374: data <= 'd0; 8375: data <= 'd0; 8376: data <= 'd0; 8377: data <= 'd0; 8378: data <= 'd0; 8379: data <= 'd0; 8380: data <= 'd0; 8381: data <= 'd0; 8382: data <= 'd0; 8383: data <= 'd0; 8384: data <= 'd0; 8385: data <= 'd0; 8386: data <= 'd0; 8387: data <= 'd0; 8388: data <= 'd0; 8389: data <= 'd0; 8390: data <= 'd0; 8391: data <= 'd0; 8392: data <= 'd0; 8393: data <= 'd0; 8394: data <= 'd0; 8395: data <= 'd0; 8396: data <= 'd0; 8397: data <= 'd0; 8398: data <= 'd0; 8399: data <= 'd0; 8400: data <= 'd0; 8401: data <= 'd0; 8402: data <= 'd0; 8403: data <= 'd0; 8404: data <= 'd0; 8405: data <= 'd0; 8406: data <= 'd0; 8407: data <= 'd0; 8408: data <= 'd0; 8409: data <= 'd0; 8410: data <= 'd0; 8411: data <= 'd0; 8412: data <= 'd0; 8413: data <= 'd0; 8414: data <= 'd0; 8415: data <= 'd0; 8416: data <= 'd0; 8417: data <= 'd0; 8418: data <= 'd0; 8419: data <= 'd0; 8420: data <= 'd0; 8421: data <= 'd0; 8422: data <= 'd0; 8423: data <= 'd0; 8424: data <= 'd0; 8425: data <= 'd0; 8426: data <= 'd0; 8427: data <= 'd0; 8428: data <= 'd0; 8429: data <= 'd0; 8430: data <= 'd0; 8431: data <= 'd0; 8432: data <= 'd0; 8433: data <= 'd0; 8434: data <= 'd0; 8435: data <= 'd0; 8436: data <= 'd0; 8437: data <= 'd0; 8438: data <= 'd0; 8439: data <= 'd0; 8440: data <= 'd0; 8441: data <= 'd0; 8442: data <= 'd0; 8443: data <= 'd0; 8444: data <= 'd0; 8445: data <= 'd0; 8446: data <= 'd0; 8447: data <= 'd0; 8448: data <= 'd0; 8449: data <= 'd0; 8450: data <= 'd0; 8451: data <= 'd0; 8452: data <= 'd0; 8453: data <= 'd0; 8454: data <= 'd0; 8455: data <= 'd0; 8456: data <= 'd0; 8457: data <= 'd0; 8458: data <= 'd0; 8459: data <= 'd1; 8460: data <= 'd1; 8461: data <= 'd1; 8462: data <= 'd1; 8463: data <= 'd0; 8464: data <= 'd0; 8465: data <= 'd0; 8466: data <= 'd0; 8467: data <= 'd0; 8468: data <= 'd0; 8469: data <= 'd0; 8470: data <= 'd0; 8471: data <= 'd0; 8472: data <= 'd0; 8473: data <= 'd0; 8474: data <= 'd0; 8475: data <= 'd0; 8476: data <= 'd0; 8477: data <= 'd0; 8478: data <= 'd0; 8479: data <= 'd0; 8480: data <= 'd0; 8481: data <= 'd0; 8482: data <= 'd0; 8483: data <= 'd0; 8484: data <= 'd0; 8485: data <= 'd0; 8486: data <= 'd0; 8487: data <= 'd0; 8488: data <= 'd0; 8489: data <= 'd0; 8490: data <= 'd0; 8491: data <= 'd0; 8492: data <= 'd0; 8493: data <= 'd0; 8494: data <= 'd0; 8495: data <= 'd0; 8496: data <= 'd0; 8497: data <= 'd0; 8498: data <= 'd0; 8499: data <= 'd0; 8500: data <= 'd0; 8501: data <= 'd0; 8502: data <= 'd0; 8503: data <= 'd0; 8504: data <= 'd0; 8505: data <= 'd0; 8506: data <= 'd0; 8507: data <= 'd0; 8508: data <= 'd0; 8509: data <= 'd0; 8510: data <= 'd0; 8511: data <= 'd0; 8512: data <= 'd0; 8513: data <= 'd0; 8514: data <= 'd0; 8515: data <= 'd0; 8516: data <= 'd0; 8517: data <= 'd0; 8518: data <= 'd0; 8519: data <= 'd0; 8520: data <= 'd0; 8521: data <= 'd0; 8522: data <= 'd0; 8523: data <= 'd0; 8524: data <= 'd0; 8525: data <= 'd0; 8526: data <= 'd0; 8527: data <= 'd0; 8528: data <= 'd0; 8529: data <= 'd0; 8530: data <= 'd0; 8531: data <= 'd0; 8532: data <= 'd0; 8533: data <= 'd0; 8534: data <= 'd0; 8535: data <= 'd0; 8536: data <= 'd0; 8537: data <= 'd0; 8538: data <= 'd0; 8539: data <= 'd0; 8540: data <= 'd0; 8541: data <= 'd0; 8542: data <= 'd0; 8543: data <= 'd0; 8544: data <= 'd0; 8545: data <= 'd0; 8546: data <= 'd0; 8547: data <= 'd0; 8548: data <= 'd0; 8549: data <= 'd0; 8550: data <= 'd0; 8551: data <= 'd0; 8552: data <= 'd0; 8553: data <= 'd0; 8554: data <= 'd0; 8555: data <= 'd0; 8556: data <= 'd0; 8557: data <= 'd0; 8558: data <= 'd0; 8559: data <= 'd0; 8560: data <= 'd0; 8561: data <= 'd0; 8562: data <= 'd0; 8563: data <= 'd0; 8564: data <= 'd0; 8565: data <= 'd0; 8566: data <= 'd0; 8567: data <= 'd0; 8568: data <= 'd0; 8569: data <= 'd0; 8570: data <= 'd0; 8571: data <= 'd0; 8572: data <= 'd0; 8573: data <= 'd0; 8574: data <= 'd0; 8575: data <= 'd0; 8576: data <= 'd0; 8577: data <= 'd0; 8578: data <= 'd0; 8579: data <= 'd0; 8580: data <= 'd0; 8581: data <= 'd0; 8582: data <= 'd0; 8583: data <= 'd0; 8584: data <= 'd0; 8585: data <= 'd0; 8586: data <= 'd0; 8587: data <= 'd0; 8588: data <= 'd1; 8589: data <= 'd1; 8590: data <= 'd0; 8591: data <= 'd0; 8592: data <= 'd0; 8593: data <= 'd0; 8594: data <= 'd0; 8595: data <= 'd0; 8596: data <= 'd0; 8597: data <= 'd0; 8598: data <= 'd0; 8599: data <= 'd0; 8600: data <= 'd0; 8601: data <= 'd0; 8602: data <= 'd0; 8603: data <= 'd0; 8604: data <= 'd0; 8605: data <= 'd0; 8606: data <= 'd0; 8607: data <= 'd0; 8608: data <= 'd0; 8609: data <= 'd0; 8610: data <= 'd0; 8611: data <= 'd0; 8612: data <= 'd0; 8613: data <= 'd0; 8614: data <= 'd0; 8615: data <= 'd0; 8616: data <= 'd0; 8617: data <= 'd0; 8618: data <= 'd0; 8619: data <= 'd0; 8620: data <= 'd0; 8621: data <= 'd0; 8622: data <= 'd0; 8623: data <= 'd0; 8624: data <= 'd0; 8625: data <= 'd0; 8626: data <= 'd0; 8627: data <= 'd0; 8628: data <= 'd0; 8629: data <= 'd0; 8630: data <= 'd0; 8631: data <= 'd0; 8632: data <= 'd0; 8633: data <= 'd0; 8634: data <= 'd0; 8635: data <= 'd0; 8636: data <= 'd0; 8637: data <= 'd0; 8638: data <= 'd0; 8639: data <= 'd0; 8640: data <= 'd0; 8641: data <= 'd0; 8642: data <= 'd0; 8643: data <= 'd0; 8644: data <= 'd0; 8645: data <= 'd0; 8646: data <= 'd0; 8647: data <= 'd0; 8648: data <= 'd0; 8649: data <= 'd0; 8650: data <= 'd0; 8651: data <= 'd0; 8652: data <= 'd0; 8653: data <= 'd0; 8654: data <= 'd0; 8655: data <= 'd0; 8656: data <= 'd0; 8657: data <= 'd0; 8658: data <= 'd0; 8659: data <= 'd0; 8660: data <= 'd0; 8661: data <= 'd0; 8662: data <= 'd0; 8663: data <= 'd0; 8664: data <= 'd0; 8665: data <= 'd0; 8666: data <= 'd0; 8667: data <= 'd0; 8668: data <= 'd0; 8669: data <= 'd0; 8670: data <= 'd0; 8671: data <= 'd0; 8672: data <= 'd0; 8673: data <= 'd0; 8674: data <= 'd0; 8675: data <= 'd0; 8676: data <= 'd0; 8677: data <= 'd0; 8678: data <= 'd0; 8679: data <= 'd0; 8680: data <= 'd0; 8681: data <= 'd0; 8682: data <= 'd0; 8683: data <= 'd0; 8684: data <= 'd0; 8685: data <= 'd0; 8686: data <= 'd0; 8687: data <= 'd0; 8688: data <= 'd0; 8689: data <= 'd0; 8690: data <= 'd0; 8691: data <= 'd0; 8692: data <= 'd0; 8693: data <= 'd0; 8694: data <= 'd0; 8695: data <= 'd0; 8696: data <= 'd0; 8697: data <= 'd0; 8698: data <= 'd0; 8699: data <= 'd0; 8700: data <= 'd0; 8701: data <= 'd0; 8702: data <= 'd0; 8703: data <= 'd0; 8704: data <= 'd0; 8705: data <= 'd0; 8706: data <= 'd0; 8707: data <= 'd0; 8708: data <= 'd0; 8709: data <= 'd0; 8710: data <= 'd0; 8711: data <= 'd0; 8712: data <= 'd0; 8713: data <= 'd0; 8714: data <= 'd0; 8715: data <= 'd0; 8716: data <= 'd1; 8717: data <= 'd0; 8718: data <= 'd0; 8719: data <= 'd0; 8720: data <= 'd0; 8721: data <= 'd0; 8722: data <= 'd0; 8723: data <= 'd0; 8724: data <= 'd0; 8725: data <= 'd0; 8726: data <= 'd0; 8727: data <= 'd0; 8728: data <= 'd0; 8729: data <= 'd0; 8730: data <= 'd0; 8731: data <= 'd0; 8732: data <= 'd0; 8733: data <= 'd0; 8734: data <= 'd0; 8735: data <= 'd0; 8736: data <= 'd0; 8737: data <= 'd0; 8738: data <= 'd0; 8739: data <= 'd0; 8740: data <= 'd0; 8741: data <= 'd0; 8742: data <= 'd0; 8743: data <= 'd0; 8744: data <= 'd0; 8745: data <= 'd0; 8746: data <= 'd0; 8747: data <= 'd0; 8748: data <= 'd0; 8749: data <= 'd0; 8750: data <= 'd0; 8751: data <= 'd0; 8752: data <= 'd0; 8753: data <= 'd0; 8754: data <= 'd0; 8755: data <= 'd0; 8756: data <= 'd0; 8757: data <= 'd0; 8758: data <= 'd0; 8759: data <= 'd0; 8760: data <= 'd0; 8761: data <= 'd0; 8762: data <= 'd0; 8763: data <= 'd0; 8764: data <= 'd0; 8765: data <= 'd0; 8766: data <= 'd0; 8767: data <= 'd0; 8768: data <= 'd0; 8769: data <= 'd0; 8770: data <= 'd0; 8771: data <= 'd0; 8772: data <= 'd0; 8773: data <= 'd0; 8774: data <= 'd0; 8775: data <= 'd0; 8776: data <= 'd0; 8777: data <= 'd0; 8778: data <= 'd0; 8779: data <= 'd0; 8780: data <= 'd0; 8781: data <= 'd0; 8782: data <= 'd0; 8783: data <= 'd0; 8784: data <= 'd0; 8785: data <= 'd0; 8786: data <= 'd0; 8787: data <= 'd0; 8788: data <= 'd0; 8789: data <= 'd0; 8790: data <= 'd0; 8791: data <= 'd0; 8792: data <= 'd0; 8793: data <= 'd0; 8794: data <= 'd0; 8795: data <= 'd0; 8796: data <= 'd0; 8797: data <= 'd0; 8798: data <= 'd0; 8799: data <= 'd0; 8800: data <= 'd0; 8801: data <= 'd0; 8802: data <= 'd0; 8803: data <= 'd0; 8804: data <= 'd0; 8805: data <= 'd0; 8806: data <= 'd0; 8807: data <= 'd0; 8808: data <= 'd0; 8809: data <= 'd0; 8810: data <= 'd0; 8811: data <= 'd0; 8812: data <= 'd0; 8813: data <= 'd0; 8814: data <= 'd0; 8815: data <= 'd0; 8816: data <= 'd0; 8817: data <= 'd0; 8818: data <= 'd0; 8819: data <= 'd0; 8820: data <= 'd0; 8821: data <= 'd0; 8822: data <= 'd0; 8823: data <= 'd0; 8824: data <= 'd0; 8825: data <= 'd0; 8826: data <= 'd0; 8827: data <= 'd0; 8828: data <= 'd0; 8829: data <= 'd0; 8830: data <= 'd0; 8831: data <= 'd0; 8832: data <= 'd0; 8833: data <= 'd0; 8834: data <= 'd0; 8835: data <= 'd0; 8836: data <= 'd0; 8837: data <= 'd0; 8838: data <= 'd0; 8839: data <= 'd0; 8840: data <= 'd0; 8841: data <= 'd0; 8842: data <= 'd0; 8843: data <= 'd1; 8844: data <= 'd1; 8845: data <= 'd0; 8846: data <= 'd0; 8847: data <= 'd0; 8848: data <= 'd0; 8849: data <= 'd0; 8850: data <= 'd0; 8851: data <= 'd0; 8852: data <= 'd0; 8853: data <= 'd0; 8854: data <= 'd0; 8855: data <= 'd0; 8856: data <= 'd0; 8857: data <= 'd0; 8858: data <= 'd0; 8859: data <= 'd0; 8860: data <= 'd0; 8861: data <= 'd0; 8862: data <= 'd0; 8863: data <= 'd0; 8864: data <= 'd0; 8865: data <= 'd0; 8866: data <= 'd0; 8867: data <= 'd0; 8868: data <= 'd0; 8869: data <= 'd0; 8870: data <= 'd0; 8871: data <= 'd0; 8872: data <= 'd0; 8873: data <= 'd0; 8874: data <= 'd0; 8875: data <= 'd0; 8876: data <= 'd0; 8877: data <= 'd0; 8878: data <= 'd0; 8879: data <= 'd0; 8880: data <= 'd0; 8881: data <= 'd0; 8882: data <= 'd0; 8883: data <= 'd0; 8884: data <= 'd0; 8885: data <= 'd0; 8886: data <= 'd0; 8887: data <= 'd0; 8888: data <= 'd0; 8889: data <= 'd0; 8890: data <= 'd0; 8891: data <= 'd0; 8892: data <= 'd0; 8893: data <= 'd0; 8894: data <= 'd0; 8895: data <= 'd0; 8896: data <= 'd0; 8897: data <= 'd0; 8898: data <= 'd0; 8899: data <= 'd0; 8900: data <= 'd0; 8901: data <= 'd0; 8902: data <= 'd0; 8903: data <= 'd0; 8904: data <= 'd0; 8905: data <= 'd0; 8906: data <= 'd0; 8907: data <= 'd0; 8908: data <= 'd0; 8909: data <= 'd0; 8910: data <= 'd0; 8911: data <= 'd0; 8912: data <= 'd0; 8913: data <= 'd0; 8914: data <= 'd0; 8915: data <= 'd0; 8916: data <= 'd0; 8917: data <= 'd0; 8918: data <= 'd0; 8919: data <= 'd0; 8920: data <= 'd0; 8921: data <= 'd0; 8922: data <= 'd0; 8923: data <= 'd0; 8924: data <= 'd0; 8925: data <= 'd0; 8926: data <= 'd0; 8927: data <= 'd0; 8928: data <= 'd0; 8929: data <= 'd0; 8930: data <= 'd0; 8931: data <= 'd0; 8932: data <= 'd0; 8933: data <= 'd0; 8934: data <= 'd0; 8935: data <= 'd0; 8936: data <= 'd0; 8937: data <= 'd0; 8938: data <= 'd0; 8939: data <= 'd0; 8940: data <= 'd0; 8941: data <= 'd0; 8942: data <= 'd0; 8943: data <= 'd0; 8944: data <= 'd0; 8945: data <= 'd0; 8946: data <= 'd0; 8947: data <= 'd0; 8948: data <= 'd0; 8949: data <= 'd0; 8950: data <= 'd0; 8951: data <= 'd0; 8952: data <= 'd0; 8953: data <= 'd0; 8954: data <= 'd0; 8955: data <= 'd0; 8956: data <= 'd0; 8957: data <= 'd0; 8958: data <= 'd0; 8959: data <= 'd0; 8960: data <= 'd0; 8961: data <= 'd0; 8962: data <= 'd0; 8963: data <= 'd0; 8964: data <= 'd0; 8965: data <= 'd0; 8966: data <= 'd0; 8967: data <= 'd0; 8968: data <= 'd0; 8969: data <= 'd0; 8970: data <= 'd0; 8971: data <= 'd1; 8972: data <= 'd0; 8973: data <= 'd0; 8974: data <= 'd0; 8975: data <= 'd0; 8976: data <= 'd0; 8977: data <= 'd0; 8978: data <= 'd0; 8979: data <= 'd0; 8980: data <= 'd0; 8981: data <= 'd0; 8982: data <= 'd0; 8983: data <= 'd0; 8984: data <= 'd0; 8985: data <= 'd0; 8986: data <= 'd0; 8987: data <= 'd0; 8988: data <= 'd0; 8989: data <= 'd0; 8990: data <= 'd0; 8991: data <= 'd0; 8992: data <= 'd0; 8993: data <= 'd0; 8994: data <= 'd0; 8995: data <= 'd0; 8996: data <= 'd0; 8997: data <= 'd0; 8998: data <= 'd0; 8999: data <= 'd0; 9000: data <= 'd0; 9001: data <= 'd0; 9002: data <= 'd0; 9003: data <= 'd0; 9004: data <= 'd0; 9005: data <= 'd0; 9006: data <= 'd0; 9007: data <= 'd0; 9008: data <= 'd0; 9009: data <= 'd0; 9010: data <= 'd0; 9011: data <= 'd0; 9012: data <= 'd0; 9013: data <= 'd0; 9014: data <= 'd0; 9015: data <= 'd0; 9016: data <= 'd0; 9017: data <= 'd0; 9018: data <= 'd0; 9019: data <= 'd0; 9020: data <= 'd0; 9021: data <= 'd0; 9022: data <= 'd0; 9023: data <= 'd0; 9024: data <= 'd0; 9025: data <= 'd0; 9026: data <= 'd0; 9027: data <= 'd0; 9028: data <= 'd0; 9029: data <= 'd0; 9030: data <= 'd0; 9031: data <= 'd0; 9032: data <= 'd0; 9033: data <= 'd0; 9034: data <= 'd0; 9035: data <= 'd0; 9036: data <= 'd0; 9037: data <= 'd0; 9038: data <= 'd0; 9039: data <= 'd0; 9040: data <= 'd0; 9041: data <= 'd0; 9042: data <= 'd0; 9043: data <= 'd0; 9044: data <= 'd0; 9045: data <= 'd0; 9046: data <= 'd0; 9047: data <= 'd0; 9048: data <= 'd0; 9049: data <= 'd0; 9050: data <= 'd0; 9051: data <= 'd0; 9052: data <= 'd0; 9053: data <= 'd0; 9054: data <= 'd0; 9055: data <= 'd0; 9056: data <= 'd0; 9057: data <= 'd0; 9058: data <= 'd0; 9059: data <= 'd0; 9060: data <= 'd0; 9061: data <= 'd0; 9062: data <= 'd0; 9063: data <= 'd0; 9064: data <= 'd0; 9065: data <= 'd0; 9066: data <= 'd0; 9067: data <= 'd0; 9068: data <= 'd0; 9069: data <= 'd0; 9070: data <= 'd0; 9071: data <= 'd0; 9072: data <= 'd0; 9073: data <= 'd0; 9074: data <= 'd0; 9075: data <= 'd0; 9076: data <= 'd0; 9077: data <= 'd0; 9078: data <= 'd0; 9079: data <= 'd0; 9080: data <= 'd0; 9081: data <= 'd0; 9082: data <= 'd0; 9083: data <= 'd0; 9084: data <= 'd0; 9085: data <= 'd0; 9086: data <= 'd0; 9087: data <= 'd0; 9088: data <= 'd0; 9089: data <= 'd0; 9090: data <= 'd0; 9091: data <= 'd0; 9092: data <= 'd0; 9093: data <= 'd0; 9094: data <= 'd0; 9095: data <= 'd0; 9096: data <= 'd0; 9097: data <= 'd0; 9098: data <= 'd0; 9099: data <= 'd1; 9100: data <= 'd0; 9101: data <= 'd0; 9102: data <= 'd0; 9103: data <= 'd0; 9104: data <= 'd0; 9105: data <= 'd0; 9106: data <= 'd0; 9107: data <= 'd0; 9108: data <= 'd0; 9109: data <= 'd0; 9110: data <= 'd0; 9111: data <= 'd0; 9112: data <= 'd0; 9113: data <= 'd0; 9114: data <= 'd0; 9115: data <= 'd0; 9116: data <= 'd0; 9117: data <= 'd0; 9118: data <= 'd0; 9119: data <= 'd0; 9120: data <= 'd0; 9121: data <= 'd0; 9122: data <= 'd0; 9123: data <= 'd0; 9124: data <= 'd0; 9125: data <= 'd0; 9126: data <= 'd0; 9127: data <= 'd0; 9128: data <= 'd0; 9129: data <= 'd0; 9130: data <= 'd0; 9131: data <= 'd0; 9132: data <= 'd0; 9133: data <= 'd0; 9134: data <= 'd0; 9135: data <= 'd0; 9136: data <= 'd0; 9137: data <= 'd0; 9138: data <= 'd0; 9139: data <= 'd0; 9140: data <= 'd0; 9141: data <= 'd0; 9142: data <= 'd0; 9143: data <= 'd0; 9144: data <= 'd0; 9145: data <= 'd0; 9146: data <= 'd0; 9147: data <= 'd0; 9148: data <= 'd0; 9149: data <= 'd0; 9150: data <= 'd0; 9151: data <= 'd0; 9152: data <= 'd0; 9153: data <= 'd0; 9154: data <= 'd0; 9155: data <= 'd0; 9156: data <= 'd0; 9157: data <= 'd0; 9158: data <= 'd0; 9159: data <= 'd0; 9160: data <= 'd0; 9161: data <= 'd0; 9162: data <= 'd0; 9163: data <= 'd0; 9164: data <= 'd0; 9165: data <= 'd0; 9166: data <= 'd0; 9167: data <= 'd0; 9168: data <= 'd0; 9169: data <= 'd0; 9170: data <= 'd0; 9171: data <= 'd0; 9172: data <= 'd0; 9173: data <= 'd0; 9174: data <= 'd0; 9175: data <= 'd0; 9176: data <= 'd0; 9177: data <= 'd0; 9178: data <= 'd0; 9179: data <= 'd0; 9180: data <= 'd0; 9181: data <= 'd0; 9182: data <= 'd0; 9183: data <= 'd0; 9184: data <= 'd0; 9185: data <= 'd0; 9186: data <= 'd0; 9187: data <= 'd0; 9188: data <= 'd0; 9189: data <= 'd0; 9190: data <= 'd0; 9191: data <= 'd0; 9192: data <= 'd0; 9193: data <= 'd0; 9194: data <= 'd0; 9195: data <= 'd0; 9196: data <= 'd0; 9197: data <= 'd0; 9198: data <= 'd0; 9199: data <= 'd0; 9200: data <= 'd0; 9201: data <= 'd0; 9202: data <= 'd0; 9203: data <= 'd0; 9204: data <= 'd0; 9205: data <= 'd0; 9206: data <= 'd0; 9207: data <= 'd0; 9208: data <= 'd0; 9209: data <= 'd0; 9210: data <= 'd0; 9211: data <= 'd0; 9212: data <= 'd0; 9213: data <= 'd0; 9214: data <= 'd0; 9215: data <= 'd0; 9216: data <= 'd0; 9217: data <= 'd0; 9218: data <= 'd0; 9219: data <= 'd0; 9220: data <= 'd0; 9221: data <= 'd0; 9222: data <= 'd0; 9223: data <= 'd0; 9224: data <= 'd0; 9225: data <= 'd0; 9226: data <= 'd0; 9227: data <= 'd1; 9228: data <= 'd0; 9229: data <= 'd0; 9230: data <= 'd0; 9231: data <= 'd0; 9232: data <= 'd0; 9233: data <= 'd0; 9234: data <= 'd0; 9235: data <= 'd0; 9236: data <= 'd0; 9237: data <= 'd0; 9238: data <= 'd0; 9239: data <= 'd0; 9240: data <= 'd0; 9241: data <= 'd0; 9242: data <= 'd0; 9243: data <= 'd0; 9244: data <= 'd0; 9245: data <= 'd0; 9246: data <= 'd0; 9247: data <= 'd0; 9248: data <= 'd0; 9249: data <= 'd0; 9250: data <= 'd0; 9251: data <= 'd0; 9252: data <= 'd0; 9253: data <= 'd0; 9254: data <= 'd0; 9255: data <= 'd0; 9256: data <= 'd0; 9257: data <= 'd0; 9258: data <= 'd0; 9259: data <= 'd0; 9260: data <= 'd0; 9261: data <= 'd0; 9262: data <= 'd0; 9263: data <= 'd0; 9264: data <= 'd0; 9265: data <= 'd0; 9266: data <= 'd0; 9267: data <= 'd0; 9268: data <= 'd0; 9269: data <= 'd0; 9270: data <= 'd0; 9271: data <= 'd0; 9272: data <= 'd0; 9273: data <= 'd0; 9274: data <= 'd0; 9275: data <= 'd0; 9276: data <= 'd0; 9277: data <= 'd0; 9278: data <= 'd0; 9279: data <= 'd0; 9280: data <= 'd0; 9281: data <= 'd0; 9282: data <= 'd0; 9283: data <= 'd0; 9284: data <= 'd0; 9285: data <= 'd0; 9286: data <= 'd0; 9287: data <= 'd0; 9288: data <= 'd0; 9289: data <= 'd0; 9290: data <= 'd0; 9291: data <= 'd0; 9292: data <= 'd0; 9293: data <= 'd0; 9294: data <= 'd0; 9295: data <= 'd0; 9296: data <= 'd0; 9297: data <= 'd0; 9298: data <= 'd0; 9299: data <= 'd0; 9300: data <= 'd0; 9301: data <= 'd0; 9302: data <= 'd0; 9303: data <= 'd0; 9304: data <= 'd0; 9305: data <= 'd0; 9306: data <= 'd0; 9307: data <= 'd0; 9308: data <= 'd0; 9309: data <= 'd0; 9310: data <= 'd0; 9311: data <= 'd0; 9312: data <= 'd0; 9313: data <= 'd0; 9314: data <= 'd0; 9315: data <= 'd0; 9316: data <= 'd0; 9317: data <= 'd0; 9318: data <= 'd0; 9319: data <= 'd0; 9320: data <= 'd0; 9321: data <= 'd0; 9322: data <= 'd0; 9323: data <= 'd0; 9324: data <= 'd0; 9325: data <= 'd0; 9326: data <= 'd0; 9327: data <= 'd0; 9328: data <= 'd0; 9329: data <= 'd0; 9330: data <= 'd0; 9331: data <= 'd0; 9332: data <= 'd0; 9333: data <= 'd0; 9334: data <= 'd0; 9335: data <= 'd0; 9336: data <= 'd0; 9337: data <= 'd0; 9338: data <= 'd0; 9339: data <= 'd0; 9340: data <= 'd0; 9341: data <= 'd0; 9342: data <= 'd0; 9343: data <= 'd0; 
default: data <= 1'bx;
        endcase
    end
assign dout = data;

endmodule