// ROMs Using Block RAM Resources.
// File: rams_sp_rom_1.v
//
module character_rom(clk, en, addr, dout);
input clk;
input en;
input [13:0] addr;
output [3:0] dout;

logic [3:0] data;

always_ff @(posedge clk) begin
    if (en)
        case(addr)
0: data <= 'd0; 1: data <= 'd0; 2: data <= 'd0; 3: data <= 'd0; 4: data <= 'd0; 5: data <= 'd0; 6: data <= 'd0; 7: data <= 'd0; 8: data <= 'd0; 9: data <= 'd0; 10: data <= 'd0; 11: data <= 'd0; 12: data <= 'd0; 13: data <= 'd0; 14: data <= 'd0; 15: data <= 'd0; 16: data <= 'd0; 17: data <= 'd0; 18: data <= 'd0; 19: data <= 'd0; 20: data <= 'd0; 21: data <= 'd0; 22: data <= 'd0; 23: data <= 'd0; 24: data <= 'd0; 25: data <= 'd0; 26: data <= 'd0; 27: data <= 'd0; 28: data <= 'd0; 29: data <= 'd0; 30: data <= 'd0; 31: data <= 'd0; 32: data <= 'd0; 33: data <= 'd0; 34: data <= 'd0; 35: data <= 'd0; 36: data <= 'd0; 37: data <= 'd0; 38: data <= 'd0; 39: data <= 'd0; 40: data <= 'd0; 41: data <= 'd0; 42: data <= 'd0; 43: data <= 'd0; 44: data <= 'd0; 45: data <= 'd0; 46: data <= 'd0; 47: data <= 'd0; 48: data <= 'd0; 49: data <= 'd0; 50: data <= 'd0; 51: data <= 'd0; 52: data <= 'd0; 53: data <= 'd0; 54: data <= 'd0; 55: data <= 'd0; 56: data <= 'd0; 57: data <= 'd0; 58: data <= 'd0; 59: data <= 'd0; 60: data <= 'd0; 61: data <= 'd0; 62: data <= 'd0; 63: data <= 'd0; 64: data <= 'd0; 65: data <= 'd0; 66: data <= 'd0; 67: data <= 'd0; 68: data <= 'd0; 69: data <= 'd0; 70: data <= 'd0; 71: data <= 'd0; 72: data <= 'd0; 73: data <= 'd0; 74: data <= 'd0; 75: data <= 'd0; 76: data <= 'd0; 77: data <= 'd0; 78: data <= 'd0; 79: data <= 'd0; 80: data <= 'd0; 81: data <= 'd0; 82: data <= 'd0; 83: data <= 'd0; 84: data <= 'd0; 85: data <= 'd0; 86: data <= 'd0; 87: data <= 'd0; 88: data <= 'd0; 89: data <= 'd0; 90: data <= 'd0; 91: data <= 'd0; 92: data <= 'd0; 93: data <= 'd0; 94: data <= 'd0; 95: data <= 'd0; 96: data <= 'd0; 97: data <= 'd0; 98: data <= 'd0; 99: data <= 'd0; 100: data <= 'd0; 101: data <= 'd0; 102: data <= 'd0; 103: data <= 'd0; 104: data <= 'd0; 105: data <= 'd0; 106: data <= 'd0; 107: data <= 'd0; 108: data <= 'd0; 109: data <= 'd0; 110: data <= 'd0; 111: data <= 'd0; 112: data <= 'd0; 113: data <= 'd0; 114: data <= 'd0; 115: data <= 'd0; 116: data <= 'd0; 117: data <= 'd0; 118: data <= 'd0; 119: data <= 'd0; 120: data <= 'd0; 121: data <= 'd0; 122: data <= 'd0; 123: data <= 'd0; 124: data <= 'd0; 125: data <= 'd0; 126: data <= 'd0; 127: data <= 'd0; 128: data <= 'd0; 129: data <= 'd0; 130: data <= 'd0; 131: data <= 'd0; 132: data <= 'd0; 133: data <= 'd0; 134: data <= 'd0; 135: data <= 'd0; 136: data <= 'd0; 137: data <= 'd0; 138: data <= 'd0; 139: data <= 'd0; 140: data <= 'd0; 141: data <= 'd0; 142: data <= 'd0; 143: data <= 'd0; 144: data <= 'd0; 145: data <= 'd0; 146: data <= 'd0; 147: data <= 'd0; 148: data <= 'd0; 149: data <= 'd0; 150: data <= 'd0; 151: data <= 'd0; 152: data <= 'd0; 153: data <= 'd0; 154: data <= 'd0; 155: data <= 'd0; 156: data <= 'd0; 157: data <= 'd0; 158: data <= 'd0; 159: data <= 'd0; 160: data <= 'd0; 161: data <= 'd0; 162: data <= 'd0; 163: data <= 'd0; 164: data <= 'd0; 165: data <= 'd0; 166: data <= 'd0; 167: data <= 'd0; 168: data <= 'd0; 169: data <= 'd0; 170: data <= 'd0; 171: data <= 'd0; 172: data <= 'd0; 173: data <= 'd0; 174: data <= 'd0; 175: data <= 'd0; 176: data <= 'd0; 177: data <= 'd0; 178: data <= 'd0; 179: data <= 'd0; 180: data <= 'd0; 181: data <= 'd0; 182: data <= 'd0; 183: data <= 'd0; 184: data <= 'd0; 185: data <= 'd0; 186: data <= 'd0; 187: data <= 'd0; 188: data <= 'd0; 189: data <= 'd0; 190: data <= 'd0; 191: data <= 'd0; 192: data <= 'd0; 193: data <= 'd0; 194: data <= 'd0; 195: data <= 'd0; 196: data <= 'd0; 197: data <= 'd0; 198: data <= 'd0; 199: data <= 'd0; 200: data <= 'd0; 201: data <= 'd0; 202: data <= 'd0; 203: data <= 'd0; 204: data <= 'd0; 205: data <= 'd0; 206: data <= 'd0; 207: data <= 'd0; 208: data <= 'd0; 209: data <= 'd0; 210: data <= 'd0; 211: data <= 'd0; 212: data <= 'd0; 213: data <= 'd0; 214: data <= 'd0; 215: data <= 'd0; 216: data <= 'd0; 217: data <= 'd0; 218: data <= 'd0; 219: data <= 'd0; 220: data <= 'd0; 221: data <= 'd0; 222: data <= 'd0; 223: data <= 'd0; 224: data <= 'd0; 225: data <= 'd0; 226: data <= 'd0; 227: data <= 'd0; 228: data <= 'd0; 229: data <= 'd0; 230: data <= 'd0; 231: data <= 'd0; 232: data <= 'd0; 233: data <= 'd0; 234: data <= 'd0; 235: data <= 'd0; 236: data <= 'd0; 237: data <= 'd0; 238: data <= 'd0; 239: data <= 'd0; 240: data <= 'd0; 241: data <= 'd0; 242: data <= 'd0; 243: data <= 'd0; 244: data <= 'd0; 245: data <= 'd0; 246: data <= 'd0; 247: data <= 'd0; 248: data <= 'd0; 249: data <= 'd0; 250: data <= 'd0; 251: data <= 'd0; 252: data <= 'd0; 253: data <= 'd0; 254: data <= 'd0; 255: data <= 'd0; 256: data <= 'd0; 257: data <= 'd0; 258: data <= 'd0; 259: data <= 'd0; 260: data <= 'd0; 261: data <= 'd0; 262: data <= 'd0; 263: data <= 'd0; 264: data <= 'd0; 265: data <= 'd0; 266: data <= 'd0; 267: data <= 'd0; 268: data <= 'd0; 269: data <= 'd0; 270: data <= 'd0; 271: data <= 'd0; 272: data <= 'd0; 273: data <= 'd0; 274: data <= 'd0; 275: data <= 'd0; 276: data <= 'd0; 277: data <= 'd0; 278: data <= 'd0; 279: data <= 'd0; 280: data <= 'd0; 281: data <= 'd0; 282: data <= 'd0; 283: data <= 'd0; 284: data <= 'd0; 285: data <= 'd0; 286: data <= 'd0; 287: data <= 'd0; 288: data <= 'd0; 289: data <= 'd0; 290: data <= 'd0; 291: data <= 'd0; 292: data <= 'd0; 293: data <= 'd0; 294: data <= 'd0; 295: data <= 'd0; 296: data <= 'd0; 297: data <= 'd0; 298: data <= 'd0; 299: data <= 'd0; 300: data <= 'd0; 301: data <= 'd2; 302: data <= 'd2; 303: data <= 'd2; 304: data <= 'd2; 305: data <= 'd2; 306: data <= 'd2; 307: data <= 'd0; 308: data <= 'd0; 309: data <= 'd0; 310: data <= 'd0; 311: data <= 'd0; 312: data <= 'd0; 313: data <= 'd0; 314: data <= 'd0; 315: data <= 'd0; 316: data <= 'd0; 317: data <= 'd0; 318: data <= 'd0; 319: data <= 'd0; 320: data <= 'd0; 321: data <= 'd0; 322: data <= 'd0; 323: data <= 'd0; 324: data <= 'd0; 325: data <= 'd0; 326: data <= 'd0; 327: data <= 'd0; 328: data <= 'd0; 329: data <= 'd0; 330: data <= 'd0; 331: data <= 'd2; 332: data <= 'd2; 333: data <= 'd6; 334: data <= 'd6; 335: data <= 'd6; 336: data <= 'd6; 337: data <= 'd6; 338: data <= 'd6; 339: data <= 'd2; 340: data <= 'd2; 341: data <= 'd0; 342: data <= 'd0; 343: data <= 'd0; 344: data <= 'd0; 345: data <= 'd0; 346: data <= 'd0; 347: data <= 'd0; 348: data <= 'd0; 349: data <= 'd0; 350: data <= 'd0; 351: data <= 'd0; 352: data <= 'd0; 353: data <= 'd0; 354: data <= 'd0; 355: data <= 'd0; 356: data <= 'd0; 357: data <= 'd0; 358: data <= 'd0; 359: data <= 'd0; 360: data <= 'd0; 361: data <= 'd0; 362: data <= 'd2; 363: data <= 'd1; 364: data <= 'd3; 365: data <= 'd6; 366: data <= 'd6; 367: data <= 'd6; 368: data <= 'd6; 369: data <= 'd6; 370: data <= 'd6; 371: data <= 'd6; 372: data <= 'd3; 373: data <= 'd2; 374: data <= 'd0; 375: data <= 'd0; 376: data <= 'd0; 377: data <= 'd0; 378: data <= 'd0; 379: data <= 'd0; 380: data <= 'd0; 381: data <= 'd0; 382: data <= 'd0; 383: data <= 'd0; 384: data <= 'd0; 385: data <= 'd0; 386: data <= 'd0; 387: data <= 'd0; 388: data <= 'd0; 389: data <= 'd0; 390: data <= 'd0; 391: data <= 'd0; 392: data <= 'd0; 393: data <= 'd2; 394: data <= 'd1; 395: data <= 'd1; 396: data <= 'd1; 397: data <= 'd3; 398: data <= 'd6; 399: data <= 'd6; 400: data <= 'd6; 401: data <= 'd6; 402: data <= 'd6; 403: data <= 'd3; 404: data <= 'd1; 405: data <= 'd1; 406: data <= 'd2; 407: data <= 'd0; 408: data <= 'd0; 409: data <= 'd0; 410: data <= 'd0; 411: data <= 'd0; 412: data <= 'd0; 413: data <= 'd0; 414: data <= 'd0; 415: data <= 'd0; 416: data <= 'd0; 417: data <= 'd0; 418: data <= 'd0; 419: data <= 'd0; 420: data <= 'd0; 421: data <= 'd0; 422: data <= 'd0; 423: data <= 'd0; 424: data <= 'd0; 425: data <= 'd2; 426: data <= 'd1; 427: data <= 'd1; 428: data <= 'd5; 429: data <= 'd5; 430: data <= 'd5; 431: data <= 'd1; 432: data <= 'd1; 433: data <= 'd1; 434: data <= 'd1; 435: data <= 'd1; 436: data <= 'd5; 437: data <= 'd5; 438: data <= 'd2; 439: data <= 'd0; 440: data <= 'd0; 441: data <= 'd0; 442: data <= 'd0; 443: data <= 'd0; 444: data <= 'd0; 445: data <= 'd0; 446: data <= 'd0; 447: data <= 'd0; 448: data <= 'd0; 449: data <= 'd0; 450: data <= 'd0; 451: data <= 'd0; 452: data <= 'd0; 453: data <= 'd0; 454: data <= 'd0; 455: data <= 'd0; 456: data <= 'd2; 457: data <= 'd1; 458: data <= 'd5; 459: data <= 'd5; 460: data <= 'd3; 461: data <= 'd6; 462: data <= 'd6; 463: data <= 'd6; 464: data <= 'd6; 465: data <= 'd6; 466: data <= 'd6; 467: data <= 'd6; 468: data <= 'd6; 469: data <= 'd3; 470: data <= 'd5; 471: data <= 'd2; 472: data <= 'd0; 473: data <= 'd0; 474: data <= 'd0; 475: data <= 'd0; 476: data <= 'd0; 477: data <= 'd0; 478: data <= 'd0; 479: data <= 'd0; 480: data <= 'd0; 481: data <= 'd0; 482: data <= 'd0; 483: data <= 'd0; 484: data <= 'd0; 485: data <= 'd0; 486: data <= 'd0; 487: data <= 'd0; 488: data <= 'd2; 489: data <= 'd5; 490: data <= 'd3; 491: data <= 'd6; 492: data <= 'd3; 493: data <= 'd1; 494: data <= 'd1; 495: data <= 'd1; 496: data <= 'd1; 497: data <= 'd1; 498: data <= 'd1; 499: data <= 'd1; 500: data <= 'd1; 501: data <= 'd1; 502: data <= 'd3; 503: data <= 'd2; 504: data <= 'd0; 505: data <= 'd0; 506: data <= 'd0; 507: data <= 'd0; 508: data <= 'd0; 509: data <= 'd0; 510: data <= 'd0; 511: data <= 'd0; 512: data <= 'd0; 513: data <= 'd0; 514: data <= 'd0; 515: data <= 'd0; 516: data <= 'd0; 517: data <= 'd0; 518: data <= 'd0; 519: data <= 'd0; 520: data <= 'd2; 521: data <= 'd5; 522: data <= 'd3; 523: data <= 'd1; 524: data <= 'd1; 525: data <= 'd1; 526: data <= 'd5; 527: data <= 'd5; 528: data <= 'd5; 529: data <= 'd5; 530: data <= 'd5; 531: data <= 'd5; 532: data <= 'd5; 533: data <= 'd1; 534: data <= 'd1; 535: data <= 'd2; 536: data <= 'd0; 537: data <= 'd0; 538: data <= 'd0; 539: data <= 'd0; 540: data <= 'd0; 541: data <= 'd0; 542: data <= 'd0; 543: data <= 'd0; 544: data <= 'd0; 545: data <= 'd0; 546: data <= 'd0; 547: data <= 'd0; 548: data <= 'd0; 549: data <= 'd0; 550: data <= 'd0; 551: data <= 'd0; 552: data <= 'd2; 553: data <= 'd6; 554: data <= 'd1; 555: data <= 'd5; 556: data <= 'd2; 557: data <= 'd2; 558: data <= 'd2; 559: data <= 'd2; 560: data <= 'd2; 561: data <= 'd2; 562: data <= 'd2; 563: data <= 'd2; 564: data <= 'd2; 565: data <= 'd2; 566: data <= 'd5; 567: data <= 'd2; 568: data <= 'd0; 569: data <= 'd0; 570: data <= 'd0; 571: data <= 'd0; 572: data <= 'd0; 573: data <= 'd0; 574: data <= 'd0; 575: data <= 'd0; 576: data <= 'd0; 577: data <= 'd0; 578: data <= 'd0; 579: data <= 'd0; 580: data <= 'd0; 581: data <= 'd0; 582: data <= 'd2; 583: data <= 'd2; 584: data <= 'd5; 585: data <= 'd6; 586: data <= 'd5; 587: data <= 'd2; 588: data <= 'd8; 589: data <= 'd8; 590: data <= 'd8; 591: data <= 'd8; 592: data <= 'd8; 593: data <= 'd9; 594: data <= 'd9; 595: data <= 'd8; 596: data <= 'd8; 597: data <= 'd8; 598: data <= 'd2; 599: data <= 'd2; 600: data <= 'd0; 601: data <= 'd0; 602: data <= 'd0; 603: data <= 'd0; 604: data <= 'd0; 605: data <= 'd0; 606: data <= 'd0; 607: data <= 'd0; 608: data <= 'd0; 609: data <= 'd0; 610: data <= 'd0; 611: data <= 'd0; 612: data <= 'd0; 613: data <= 'd0; 614: data <= 'd2; 615: data <= 'd3; 616: data <= 'd6; 617: data <= 'd3; 618: data <= 'd2; 619: data <= 'd8; 620: data <= 'd8; 621: data <= 'd9; 622: data <= 'd9; 623: data <= 'd10; 624: data <= 'd2; 625: data <= 'd9; 626: data <= 'd11; 627: data <= 'd10; 628: data <= 'd2; 629: data <= 'd9; 630: data <= 'd2; 631: data <= 'd2; 632: data <= 'd0; 633: data <= 'd0; 634: data <= 'd0; 635: data <= 'd0; 636: data <= 'd0; 637: data <= 'd0; 638: data <= 'd0; 639: data <= 'd0; 640: data <= 'd0; 641: data <= 'd0; 642: data <= 'd0; 643: data <= 'd0; 644: data <= 'd0; 645: data <= 'd0; 646: data <= 'd2; 647: data <= 'd1; 648: data <= 'd3; 649: data <= 'd1; 650: data <= 'd2; 651: data <= 'd10; 652: data <= 'd10; 653: data <= 'd9; 654: data <= 'd10; 655: data <= 'd10; 656: data <= 'd11; 657: data <= 'd10; 658: data <= 'd11; 659: data <= 'd11; 660: data <= 'd10; 661: data <= 'd10; 662: data <= 'd2; 663: data <= 'd0; 664: data <= 'd0; 665: data <= 'd0; 666: data <= 'd0; 667: data <= 'd0; 668: data <= 'd0; 669: data <= 'd0; 670: data <= 'd0; 671: data <= 'd0; 672: data <= 'd0; 673: data <= 'd0; 674: data <= 'd0; 675: data <= 'd0; 676: data <= 'd0; 677: data <= 'd0; 678: data <= 'd0; 679: data <= 'd2; 680: data <= 'd1; 681: data <= 'd5; 682: data <= 'd2; 683: data <= 'd8; 684: data <= 'd9; 685: data <= 'd9; 686: data <= 'd10; 687: data <= 'd10; 688: data <= 'd10; 689: data <= 'd10; 690: data <= 'd8; 691: data <= 'd8; 692: data <= 'd10; 693: data <= 'd9; 694: data <= 'd2; 695: data <= 'd0; 696: data <= 'd0; 697: data <= 'd0; 698: data <= 'd0; 699: data <= 'd0; 700: data <= 'd0; 701: data <= 'd0; 702: data <= 'd0; 703: data <= 'd0; 704: data <= 'd0; 705: data <= 'd0; 706: data <= 'd0; 707: data <= 'd0; 708: data <= 'd0; 709: data <= 'd0; 710: data <= 'd0; 711: data <= 'd0; 712: data <= 'd2; 713: data <= 'd2; 714: data <= 'd2; 715: data <= 'd8; 716: data <= 'd8; 717: data <= 'd9; 718: data <= 'd9; 719: data <= 'd10; 720: data <= 'd10; 721: data <= 'd10; 722: data <= 'd9; 723: data <= 'd9; 724: data <= 'd10; 725: data <= 'd9; 726: data <= 'd2; 727: data <= 'd0; 728: data <= 'd0; 729: data <= 'd0; 730: data <= 'd0; 731: data <= 'd0; 732: data <= 'd0; 733: data <= 'd0; 734: data <= 'd0; 735: data <= 'd0; 736: data <= 'd0; 737: data <= 'd0; 738: data <= 'd0; 739: data <= 'd0; 740: data <= 'd0; 741: data <= 'd0; 742: data <= 'd0; 743: data <= 'd0; 744: data <= 'd0; 745: data <= 'd0; 746: data <= 'd0; 747: data <= 'd2; 748: data <= 'd5; 749: data <= 'd5; 750: data <= 'd8; 751: data <= 'd9; 752: data <= 'd9; 753: data <= 'd9; 754: data <= 'd9; 755: data <= 'd9; 756: data <= 'd9; 757: data <= 'd2; 758: data <= 'd0; 759: data <= 'd0; 760: data <= 'd0; 761: data <= 'd0; 762: data <= 'd0; 763: data <= 'd0; 764: data <= 'd0; 765: data <= 'd0; 766: data <= 'd0; 767: data <= 'd0; 768: data <= 'd0; 769: data <= 'd0; 770: data <= 'd0; 771: data <= 'd0; 772: data <= 'd0; 773: data <= 'd0; 774: data <= 'd0; 775: data <= 'd0; 776: data <= 'd0; 777: data <= 'd0; 778: data <= 'd2; 779: data <= 'd7; 780: data <= 'd1; 781: data <= 'd1; 782: data <= 'd1; 783: data <= 'd3; 784: data <= 'd3; 785: data <= 'd3; 786: data <= 'd5; 787: data <= 'd5; 788: data <= 'd3; 789: data <= 'd1; 790: data <= 'd2; 791: data <= 'd0; 792: data <= 'd0; 793: data <= 'd0; 794: data <= 'd0; 795: data <= 'd0; 796: data <= 'd0; 797: data <= 'd0; 798: data <= 'd0; 799: data <= 'd0; 800: data <= 'd0; 801: data <= 'd0; 802: data <= 'd0; 803: data <= 'd0; 804: data <= 'd0; 805: data <= 'd0; 806: data <= 'd0; 807: data <= 'd0; 808: data <= 'd0; 809: data <= 'd0; 810: data <= 'd2; 811: data <= 'd7; 812: data <= 'd7; 813: data <= 'd1; 814: data <= 'd1; 815: data <= 'd3; 816: data <= 'd3; 817: data <= 'd3; 818: data <= 'd1; 819: data <= 'd1; 820: data <= 'd3; 821: data <= 'd1; 822: data <= 'd2; 823: data <= 'd0; 824: data <= 'd0; 825: data <= 'd0; 826: data <= 'd0; 827: data <= 'd0; 828: data <= 'd0; 829: data <= 'd0; 830: data <= 'd0; 831: data <= 'd0; 832: data <= 'd0; 833: data <= 'd0; 834: data <= 'd0; 835: data <= 'd0; 836: data <= 'd0; 837: data <= 'd0; 838: data <= 'd0; 839: data <= 'd0; 840: data <= 'd0; 841: data <= 'd2; 842: data <= 'd9; 843: data <= 'd9; 844: data <= 'd7; 845: data <= 'd1; 846: data <= 'd1; 847: data <= 'd1; 848: data <= 'd3; 849: data <= 'd3; 850: data <= 'd1; 851: data <= 'd1; 852: data <= 'd1; 853: data <= 'd1; 854: data <= 'd8; 855: data <= 'd2; 856: data <= 'd0; 857: data <= 'd0; 858: data <= 'd0; 859: data <= 'd0; 860: data <= 'd0; 861: data <= 'd0; 862: data <= 'd0; 863: data <= 'd0; 864: data <= 'd0; 865: data <= 'd0; 866: data <= 'd0; 867: data <= 'd0; 868: data <= 'd0; 869: data <= 'd0; 870: data <= 'd0; 871: data <= 'd0; 872: data <= 'd0; 873: data <= 'd2; 874: data <= 'd9; 875: data <= 'd9; 876: data <= 'd2; 877: data <= 'd2; 878: data <= 'd2; 879: data <= 'd2; 880: data <= 'd2; 881: data <= 'd5; 882: data <= 'd5; 883: data <= 'd5; 884: data <= 'd2; 885: data <= 'd2; 886: data <= 'd8; 887: data <= 'd2; 888: data <= 'd0; 889: data <= 'd0; 890: data <= 'd0; 891: data <= 'd0; 892: data <= 'd0; 893: data <= 'd0; 894: data <= 'd0; 895: data <= 'd0; 896: data <= 'd0; 897: data <= 'd0; 898: data <= 'd0; 899: data <= 'd0; 900: data <= 'd0; 901: data <= 'd0; 902: data <= 'd0; 903: data <= 'd0; 904: data <= 'd0; 905: data <= 'd0; 906: data <= 'd2; 907: data <= 'd2; 908: data <= 'd2; 909: data <= 'd1; 910: data <= 'd1; 911: data <= 'd3; 912: data <= 'd3; 913: data <= 'd3; 914: data <= 'd3; 915: data <= 'd3; 916: data <= 'd3; 917: data <= 'd2; 918: data <= 'd2; 919: data <= 'd0; 920: data <= 'd0; 921: data <= 'd0; 922: data <= 'd0; 923: data <= 'd0; 924: data <= 'd0; 925: data <= 'd0; 926: data <= 'd0; 927: data <= 'd0; 928: data <= 'd0; 929: data <= 'd0; 930: data <= 'd0; 931: data <= 'd0; 932: data <= 'd0; 933: data <= 'd0; 934: data <= 'd0; 935: data <= 'd0; 936: data <= 'd0; 937: data <= 'd0; 938: data <= 'd0; 939: data <= 'd0; 940: data <= 'd2; 941: data <= 'd4; 942: data <= 'd7; 943: data <= 'd7; 944: data <= 'd2; 945: data <= 'd2; 946: data <= 'd5; 947: data <= 'd5; 948: data <= 'd4; 949: data <= 'd2; 950: data <= 'd0; 951: data <= 'd0; 952: data <= 'd0; 953: data <= 'd0; 954: data <= 'd0; 955: data <= 'd0; 956: data <= 'd0; 957: data <= 'd0; 958: data <= 'd0; 959: data <= 'd0; 960: data <= 'd0; 961: data <= 'd0; 962: data <= 'd0; 963: data <= 'd0; 964: data <= 'd0; 965: data <= 'd0; 966: data <= 'd0; 967: data <= 'd0; 968: data <= 'd0; 969: data <= 'd0; 970: data <= 'd0; 971: data <= 'd0; 972: data <= 'd2; 973: data <= 'd4; 974: data <= 'd7; 975: data <= 'd2; 976: data <= 'd0; 977: data <= 'd0; 978: data <= 'd2; 979: data <= 'd4; 980: data <= 'd4; 981: data <= 'd2; 982: data <= 'd0; 983: data <= 'd0; 984: data <= 'd0; 985: data <= 'd0; 986: data <= 'd0; 987: data <= 'd0; 988: data <= 'd0; 989: data <= 'd0; 990: data <= 'd0; 991: data <= 'd0; 992: data <= 'd0; 993: data <= 'd0; 994: data <= 'd0; 995: data <= 'd0; 996: data <= 'd0; 997: data <= 'd0; 998: data <= 'd0; 999: data <= 'd0; 1000: data <= 'd0; 1001: data <= 'd0; 1002: data <= 'd0; 1003: data <= 'd0; 1004: data <= 'd2; 1005: data <= 'd2; 1006: data <= 'd2; 1007: data <= 'd0; 1008: data <= 'd0; 1009: data <= 'd0; 1010: data <= 'd2; 1011: data <= 'd2; 1012: data <= 'd2; 1013: data <= 'd0; 1014: data <= 'd0; 1015: data <= 'd0; 1016: data <= 'd0; 1017: data <= 'd0; 1018: data <= 'd0; 1019: data <= 'd0; 1020: data <= 'd0; 1021: data <= 'd0; 1022: data <= 'd0; 1023: data <= 'd0; 1024: data <= 'd0; 1025: data <= 'd0; 1026: data <= 'd0; 1027: data <= 'd0; 1028: data <= 'd0; 1029: data <= 'd0; 1030: data <= 'd0; 1031: data <= 'd0; 1032: data <= 'd0; 1033: data <= 'd0; 1034: data <= 'd0; 1035: data <= 'd0; 1036: data <= 'd0; 1037: data <= 'd0; 1038: data <= 'd0; 1039: data <= 'd0; 1040: data <= 'd0; 1041: data <= 'd0; 1042: data <= 'd0; 1043: data <= 'd0; 1044: data <= 'd0; 1045: data <= 'd0; 1046: data <= 'd0; 1047: data <= 'd0; 1048: data <= 'd0; 1049: data <= 'd0; 1050: data <= 'd0; 1051: data <= 'd0; 1052: data <= 'd0; 1053: data <= 'd0; 1054: data <= 'd0; 1055: data <= 'd0; 1056: data <= 'd0; 1057: data <= 'd0; 1058: data <= 'd0; 1059: data <= 'd0; 1060: data <= 'd0; 1061: data <= 'd0; 1062: data <= 'd0; 1063: data <= 'd0; 1064: data <= 'd0; 1065: data <= 'd0; 1066: data <= 'd0; 1067: data <= 'd0; 1068: data <= 'd0; 1069: data <= 'd0; 1070: data <= 'd0; 1071: data <= 'd0; 1072: data <= 'd0; 1073: data <= 'd0; 1074: data <= 'd0; 1075: data <= 'd0; 1076: data <= 'd0; 1077: data <= 'd0; 1078: data <= 'd0; 1079: data <= 'd0; 1080: data <= 'd0; 1081: data <= 'd0; 1082: data <= 'd0; 1083: data <= 'd0; 1084: data <= 'd0; 1085: data <= 'd0; 1086: data <= 'd0; 1087: data <= 'd0; 1088: data <= 'd0; 1089: data <= 'd0; 1090: data <= 'd0; 1091: data <= 'd0; 1092: data <= 'd0; 1093: data <= 'd0; 1094: data <= 'd0; 1095: data <= 'd0; 1096: data <= 'd0; 1097: data <= 'd0; 1098: data <= 'd0; 1099: data <= 'd0; 1100: data <= 'd0; 1101: data <= 'd0; 1102: data <= 'd0; 1103: data <= 'd0; 1104: data <= 'd0; 1105: data <= 'd0; 1106: data <= 'd0; 1107: data <= 'd0; 1108: data <= 'd0; 1109: data <= 'd0; 1110: data <= 'd0; 1111: data <= 'd0; 1112: data <= 'd0; 1113: data <= 'd0; 1114: data <= 'd0; 1115: data <= 'd0; 1116: data <= 'd0; 1117: data <= 'd0; 1118: data <= 'd0; 1119: data <= 'd0; 1120: data <= 'd0; 1121: data <= 'd0; 1122: data <= 'd0; 1123: data <= 'd0; 1124: data <= 'd0; 1125: data <= 'd0; 1126: data <= 'd0; 1127: data <= 'd0; 1128: data <= 'd0; 1129: data <= 'd0; 1130: data <= 'd0; 1131: data <= 'd0; 1132: data <= 'd0; 1133: data <= 'd0; 1134: data <= 'd0; 1135: data <= 'd0; 1136: data <= 'd0; 1137: data <= 'd0; 1138: data <= 'd0; 1139: data <= 'd0; 1140: data <= 'd0; 1141: data <= 'd0; 1142: data <= 'd0; 1143: data <= 'd0; 1144: data <= 'd0; 1145: data <= 'd0; 1146: data <= 'd0; 1147: data <= 'd0; 1148: data <= 'd0; 1149: data <= 'd0; 1150: data <= 'd0; 1151: data <= 'd0; 1152: data <= 'd0; 1153: data <= 'd0; 1154: data <= 'd0; 1155: data <= 'd0; 1156: data <= 'd0; 1157: data <= 'd0; 1158: data <= 'd0; 1159: data <= 'd0; 1160: data <= 'd0; 1161: data <= 'd0; 1162: data <= 'd0; 1163: data <= 'd0; 1164: data <= 'd0; 1165: data <= 'd0; 1166: data <= 'd0; 1167: data <= 'd0; 1168: data <= 'd0; 1169: data <= 'd0; 1170: data <= 'd0; 1171: data <= 'd0; 1172: data <= 'd0; 1173: data <= 'd0; 1174: data <= 'd0; 1175: data <= 'd0; 1176: data <= 'd0; 1177: data <= 'd0; 1178: data <= 'd0; 1179: data <= 'd0; 1180: data <= 'd0; 1181: data <= 'd0; 1182: data <= 'd0; 1183: data <= 'd0; 1184: data <= 'd0; 1185: data <= 'd0; 1186: data <= 'd0; 1187: data <= 'd0; 1188: data <= 'd0; 1189: data <= 'd0; 1190: data <= 'd0; 1191: data <= 'd0; 1192: data <= 'd0; 1193: data <= 'd0; 1194: data <= 'd0; 1195: data <= 'd0; 1196: data <= 'd0; 1197: data <= 'd0; 1198: data <= 'd0; 1199: data <= 'd0; 1200: data <= 'd0; 1201: data <= 'd0; 1202: data <= 'd0; 1203: data <= 'd0; 1204: data <= 'd0; 1205: data <= 'd0; 1206: data <= 'd0; 1207: data <= 'd0; 1208: data <= 'd0; 1209: data <= 'd0; 1210: data <= 'd0; 1211: data <= 'd0; 1212: data <= 'd0; 1213: data <= 'd0; 1214: data <= 'd0; 1215: data <= 'd0; 1216: data <= 'd0; 1217: data <= 'd0; 1218: data <= 'd0; 1219: data <= 'd0; 1220: data <= 'd0; 1221: data <= 'd0; 1222: data <= 'd0; 1223: data <= 'd0; 1224: data <= 'd0; 1225: data <= 'd0; 1226: data <= 'd0; 1227: data <= 'd0; 1228: data <= 'd0; 1229: data <= 'd0; 1230: data <= 'd0; 1231: data <= 'd0; 1232: data <= 'd0; 1233: data <= 'd0; 1234: data <= 'd0; 1235: data <= 'd0; 1236: data <= 'd0; 1237: data <= 'd0; 1238: data <= 'd0; 1239: data <= 'd0; 1240: data <= 'd0; 1241: data <= 'd0; 1242: data <= 'd0; 1243: data <= 'd0; 1244: data <= 'd0; 1245: data <= 'd0; 1246: data <= 'd0; 1247: data <= 'd0; 1248: data <= 'd0; 1249: data <= 'd0; 1250: data <= 'd0; 1251: data <= 'd0; 1252: data <= 'd0; 1253: data <= 'd0; 1254: data <= 'd0; 1255: data <= 'd0; 1256: data <= 'd0; 1257: data <= 'd0; 1258: data <= 'd0; 1259: data <= 'd0; 1260: data <= 'd0; 1261: data <= 'd0; 1262: data <= 'd0; 1263: data <= 'd0; 1264: data <= 'd0; 1265: data <= 'd0; 1266: data <= 'd0; 1267: data <= 'd0; 1268: data <= 'd0; 1269: data <= 'd0; 1270: data <= 'd0; 1271: data <= 'd0; 1272: data <= 'd0; 1273: data <= 'd0; 1274: data <= 'd0; 1275: data <= 'd0; 1276: data <= 'd0; 1277: data <= 'd0; 1278: data <= 'd0; 1279: data <= 'd0; 1280: data <= 'd0; 1281: data <= 'd0; 1282: data <= 'd0; 1283: data <= 'd0; 1284: data <= 'd0; 1285: data <= 'd0; 1286: data <= 'd0; 1287: data <= 'd0; 1288: data <= 'd0; 1289: data <= 'd0; 1290: data <= 'd0; 1291: data <= 'd0; 1292: data <= 'd0; 1293: data <= 'd2; 1294: data <= 'd2; 1295: data <= 'd2; 1296: data <= 'd2; 1297: data <= 'd2; 1298: data <= 'd2; 1299: data <= 'd0; 1300: data <= 'd0; 1301: data <= 'd0; 1302: data <= 'd0; 1303: data <= 'd0; 1304: data <= 'd0; 1305: data <= 'd0; 1306: data <= 'd0; 1307: data <= 'd0; 1308: data <= 'd0; 1309: data <= 'd0; 1310: data <= 'd0; 1311: data <= 'd0; 1312: data <= 'd0; 1313: data <= 'd0; 1314: data <= 'd0; 1315: data <= 'd0; 1316: data <= 'd0; 1317: data <= 'd0; 1318: data <= 'd0; 1319: data <= 'd0; 1320: data <= 'd0; 1321: data <= 'd0; 1322: data <= 'd0; 1323: data <= 'd2; 1324: data <= 'd2; 1325: data <= 'd6; 1326: data <= 'd6; 1327: data <= 'd6; 1328: data <= 'd6; 1329: data <= 'd6; 1330: data <= 'd6; 1331: data <= 'd2; 1332: data <= 'd2; 1333: data <= 'd0; 1334: data <= 'd0; 1335: data <= 'd0; 1336: data <= 'd0; 1337: data <= 'd0; 1338: data <= 'd0; 1339: data <= 'd0; 1340: data <= 'd0; 1341: data <= 'd0; 1342: data <= 'd0; 1343: data <= 'd0; 1344: data <= 'd0; 1345: data <= 'd0; 1346: data <= 'd0; 1347: data <= 'd0; 1348: data <= 'd0; 1349: data <= 'd0; 1350: data <= 'd0; 1351: data <= 'd0; 1352: data <= 'd0; 1353: data <= 'd0; 1354: data <= 'd2; 1355: data <= 'd1; 1356: data <= 'd3; 1357: data <= 'd6; 1358: data <= 'd6; 1359: data <= 'd6; 1360: data <= 'd6; 1361: data <= 'd6; 1362: data <= 'd6; 1363: data <= 'd6; 1364: data <= 'd3; 1365: data <= 'd2; 1366: data <= 'd0; 1367: data <= 'd0; 1368: data <= 'd0; 1369: data <= 'd0; 1370: data <= 'd0; 1371: data <= 'd0; 1372: data <= 'd0; 1373: data <= 'd0; 1374: data <= 'd0; 1375: data <= 'd0; 1376: data <= 'd0; 1377: data <= 'd0; 1378: data <= 'd0; 1379: data <= 'd0; 1380: data <= 'd0; 1381: data <= 'd0; 1382: data <= 'd0; 1383: data <= 'd0; 1384: data <= 'd0; 1385: data <= 'd2; 1386: data <= 'd1; 1387: data <= 'd1; 1388: data <= 'd1; 1389: data <= 'd3; 1390: data <= 'd6; 1391: data <= 'd6; 1392: data <= 'd6; 1393: data <= 'd6; 1394: data <= 'd6; 1395: data <= 'd3; 1396: data <= 'd1; 1397: data <= 'd1; 1398: data <= 'd2; 1399: data <= 'd0; 1400: data <= 'd0; 1401: data <= 'd0; 1402: data <= 'd0; 1403: data <= 'd0; 1404: data <= 'd0; 1405: data <= 'd0; 1406: data <= 'd0; 1407: data <= 'd0; 1408: data <= 'd0; 1409: data <= 'd0; 1410: data <= 'd0; 1411: data <= 'd0; 1412: data <= 'd0; 1413: data <= 'd0; 1414: data <= 'd0; 1415: data <= 'd0; 1416: data <= 'd0; 1417: data <= 'd2; 1418: data <= 'd1; 1419: data <= 'd1; 1420: data <= 'd5; 1421: data <= 'd5; 1422: data <= 'd5; 1423: data <= 'd1; 1424: data <= 'd1; 1425: data <= 'd1; 1426: data <= 'd1; 1427: data <= 'd1; 1428: data <= 'd5; 1429: data <= 'd5; 1430: data <= 'd2; 1431: data <= 'd0; 1432: data <= 'd0; 1433: data <= 'd0; 1434: data <= 'd0; 1435: data <= 'd0; 1436: data <= 'd0; 1437: data <= 'd0; 1438: data <= 'd0; 1439: data <= 'd0; 1440: data <= 'd0; 1441: data <= 'd0; 1442: data <= 'd0; 1443: data <= 'd0; 1444: data <= 'd0; 1445: data <= 'd0; 1446: data <= 'd0; 1447: data <= 'd0; 1448: data <= 'd2; 1449: data <= 'd1; 1450: data <= 'd5; 1451: data <= 'd5; 1452: data <= 'd3; 1453: data <= 'd6; 1454: data <= 'd6; 1455: data <= 'd6; 1456: data <= 'd6; 1457: data <= 'd6; 1458: data <= 'd6; 1459: data <= 'd6; 1460: data <= 'd6; 1461: data <= 'd3; 1462: data <= 'd5; 1463: data <= 'd2; 1464: data <= 'd0; 1465: data <= 'd0; 1466: data <= 'd0; 1467: data <= 'd0; 1468: data <= 'd0; 1469: data <= 'd0; 1470: data <= 'd0; 1471: data <= 'd0; 1472: data <= 'd0; 1473: data <= 'd0; 1474: data <= 'd0; 1475: data <= 'd0; 1476: data <= 'd0; 1477: data <= 'd0; 1478: data <= 'd0; 1479: data <= 'd0; 1480: data <= 'd2; 1481: data <= 'd5; 1482: data <= 'd3; 1483: data <= 'd6; 1484: data <= 'd3; 1485: data <= 'd1; 1486: data <= 'd1; 1487: data <= 'd1; 1488: data <= 'd1; 1489: data <= 'd1; 1490: data <= 'd1; 1491: data <= 'd1; 1492: data <= 'd1; 1493: data <= 'd1; 1494: data <= 'd3; 1495: data <= 'd2; 1496: data <= 'd0; 1497: data <= 'd0; 1498: data <= 'd0; 1499: data <= 'd0; 1500: data <= 'd0; 1501: data <= 'd0; 1502: data <= 'd0; 1503: data <= 'd0; 1504: data <= 'd0; 1505: data <= 'd0; 1506: data <= 'd0; 1507: data <= 'd0; 1508: data <= 'd0; 1509: data <= 'd0; 1510: data <= 'd0; 1511: data <= 'd0; 1512: data <= 'd2; 1513: data <= 'd5; 1514: data <= 'd3; 1515: data <= 'd1; 1516: data <= 'd1; 1517: data <= 'd1; 1518: data <= 'd5; 1519: data <= 'd5; 1520: data <= 'd5; 1521: data <= 'd5; 1522: data <= 'd5; 1523: data <= 'd5; 1524: data <= 'd5; 1525: data <= 'd1; 1526: data <= 'd1; 1527: data <= 'd2; 1528: data <= 'd0; 1529: data <= 'd0; 1530: data <= 'd0; 1531: data <= 'd0; 1532: data <= 'd0; 1533: data <= 'd0; 1534: data <= 'd0; 1535: data <= 'd0; 1536: data <= 'd0; 1537: data <= 'd0; 1538: data <= 'd0; 1539: data <= 'd0; 1540: data <= 'd0; 1541: data <= 'd0; 1542: data <= 'd0; 1543: data <= 'd0; 1544: data <= 'd2; 1545: data <= 'd6; 1546: data <= 'd1; 1547: data <= 'd5; 1548: data <= 'd2; 1549: data <= 'd2; 1550: data <= 'd2; 1551: data <= 'd2; 1552: data <= 'd2; 1553: data <= 'd2; 1554: data <= 'd2; 1555: data <= 'd2; 1556: data <= 'd2; 1557: data <= 'd2; 1558: data <= 'd5; 1559: data <= 'd2; 1560: data <= 'd0; 1561: data <= 'd0; 1562: data <= 'd0; 1563: data <= 'd0; 1564: data <= 'd0; 1565: data <= 'd0; 1566: data <= 'd0; 1567: data <= 'd0; 1568: data <= 'd0; 1569: data <= 'd0; 1570: data <= 'd0; 1571: data <= 'd0; 1572: data <= 'd0; 1573: data <= 'd0; 1574: data <= 'd2; 1575: data <= 'd2; 1576: data <= 'd2; 1577: data <= 'd1; 1578: data <= 'd5; 1579: data <= 'd2; 1580: data <= 'd8; 1581: data <= 'd8; 1582: data <= 'd8; 1583: data <= 'd8; 1584: data <= 'd8; 1585: data <= 'd9; 1586: data <= 'd9; 1587: data <= 'd8; 1588: data <= 'd8; 1589: data <= 'd8; 1590: data <= 'd2; 1591: data <= 'd2; 1592: data <= 'd0; 1593: data <= 'd0; 1594: data <= 'd0; 1595: data <= 'd0; 1596: data <= 'd0; 1597: data <= 'd0; 1598: data <= 'd0; 1599: data <= 'd0; 1600: data <= 'd0; 1601: data <= 'd0; 1602: data <= 'd0; 1603: data <= 'd0; 1604: data <= 'd0; 1605: data <= 'd0; 1606: data <= 'd2; 1607: data <= 'd1; 1608: data <= 'd2; 1609: data <= 'd1; 1610: data <= 'd2; 1611: data <= 'd8; 1612: data <= 'd8; 1613: data <= 'd9; 1614: data <= 'd9; 1615: data <= 'd2; 1616: data <= 'd9; 1617: data <= 'd11; 1618: data <= 'd11; 1619: data <= 'd10; 1620: data <= 'd2; 1621: data <= 'd9; 1622: data <= 'd2; 1623: data <= 'd2; 1624: data <= 'd0; 1625: data <= 'd0; 1626: data <= 'd0; 1627: data <= 'd0; 1628: data <= 'd0; 1629: data <= 'd0; 1630: data <= 'd0; 1631: data <= 'd0; 1632: data <= 'd0; 1633: data <= 'd0; 1634: data <= 'd0; 1635: data <= 'd0; 1636: data <= 'd0; 1637: data <= 'd0; 1638: data <= 'd2; 1639: data <= 'd5; 1640: data <= 'd1; 1641: data <= 'd2; 1642: data <= 'd9; 1643: data <= 'd10; 1644: data <= 'd9; 1645: data <= 'd9; 1646: data <= 'd10; 1647: data <= 'd11; 1648: data <= 'd10; 1649: data <= 'd11; 1650: data <= 'd11; 1651: data <= 'd10; 1652: data <= 'd11; 1653: data <= 'd10; 1654: data <= 'd9; 1655: data <= 'd2; 1656: data <= 'd0; 1657: data <= 'd0; 1658: data <= 'd0; 1659: data <= 'd0; 1660: data <= 'd0; 1661: data <= 'd0; 1662: data <= 'd0; 1663: data <= 'd0; 1664: data <= 'd0; 1665: data <= 'd0; 1666: data <= 'd0; 1667: data <= 'd0; 1668: data <= 'd0; 1669: data <= 'd0; 1670: data <= 'd0; 1671: data <= 'd2; 1672: data <= 'd5; 1673: data <= 'd5; 1674: data <= 'd2; 1675: data <= 'd8; 1676: data <= 'd9; 1677: data <= 'd9; 1678: data <= 'd10; 1679: data <= 'd10; 1680: data <= 'd10; 1681: data <= 'd8; 1682: data <= 'd8; 1683: data <= 'd10; 1684: data <= 'd10; 1685: data <= 'd9; 1686: data <= 'd2; 1687: data <= 'd0; 1688: data <= 'd0; 1689: data <= 'd0; 1690: data <= 'd0; 1691: data <= 'd0; 1692: data <= 'd0; 1693: data <= 'd0; 1694: data <= 'd0; 1695: data <= 'd0; 1696: data <= 'd0; 1697: data <= 'd0; 1698: data <= 'd0; 1699: data <= 'd0; 1700: data <= 'd0; 1701: data <= 'd0; 1702: data <= 'd0; 1703: data <= 'd0; 1704: data <= 'd2; 1705: data <= 'd2; 1706: data <= 'd2; 1707: data <= 'd8; 1708: data <= 'd8; 1709: data <= 'd9; 1710: data <= 'd9; 1711: data <= 'd10; 1712: data <= 'd10; 1713: data <= 'd9; 1714: data <= 'd9; 1715: data <= 'd10; 1716: data <= 'd10; 1717: data <= 'd9; 1718: data <= 'd2; 1719: data <= 'd0; 1720: data <= 'd0; 1721: data <= 'd0; 1722: data <= 'd0; 1723: data <= 'd0; 1724: data <= 'd0; 1725: data <= 'd0; 1726: data <= 'd0; 1727: data <= 'd0; 1728: data <= 'd0; 1729: data <= 'd0; 1730: data <= 'd0; 1731: data <= 'd0; 1732: data <= 'd0; 1733: data <= 'd0; 1734: data <= 'd0; 1735: data <= 'd0; 1736: data <= 'd0; 1737: data <= 'd0; 1738: data <= 'd2; 1739: data <= 'd2; 1740: data <= 'd5; 1741: data <= 'd5; 1742: data <= 'd8; 1743: data <= 'd9; 1744: data <= 'd9; 1745: data <= 'd9; 1746: data <= 'd9; 1747: data <= 'd9; 1748: data <= 'd9; 1749: data <= 'd5; 1750: data <= 'd2; 1751: data <= 'd0; 1752: data <= 'd0; 1753: data <= 'd0; 1754: data <= 'd0; 1755: data <= 'd0; 1756: data <= 'd0; 1757: data <= 'd0; 1758: data <= 'd0; 1759: data <= 'd0; 1760: data <= 'd0; 1761: data <= 'd0; 1762: data <= 'd0; 1763: data <= 'd0; 1764: data <= 'd0; 1765: data <= 'd0; 1766: data <= 'd0; 1767: data <= 'd0; 1768: data <= 'd0; 1769: data <= 'd2; 1770: data <= 'd7; 1771: data <= 'd1; 1772: data <= 'd1; 1773: data <= 'd1; 1774: data <= 'd3; 1775: data <= 'd3; 1776: data <= 'd3; 1777: data <= 'd5; 1778: data <= 'd5; 1779: data <= 'd3; 1780: data <= 'd3; 1781: data <= 'd1; 1782: data <= 'd2; 1783: data <= 'd0; 1784: data <= 'd0; 1785: data <= 'd0; 1786: data <= 'd0; 1787: data <= 'd0; 1788: data <= 'd0; 1789: data <= 'd0; 1790: data <= 'd0; 1791: data <= 'd0; 1792: data <= 'd0; 1793: data <= 'd0; 1794: data <= 'd0; 1795: data <= 'd0; 1796: data <= 'd0; 1797: data <= 'd0; 1798: data <= 'd0; 1799: data <= 'd0; 1800: data <= 'd0; 1801: data <= 'd2; 1802: data <= 'd7; 1803: data <= 'd7; 1804: data <= 'd5; 1805: data <= 'd1; 1806: data <= 'd3; 1807: data <= 'd3; 1808: data <= 'd3; 1809: data <= 'd1; 1810: data <= 'd1; 1811: data <= 'd3; 1812: data <= 'd3; 1813: data <= 'd1; 1814: data <= 'd2; 1815: data <= 'd0; 1816: data <= 'd0; 1817: data <= 'd0; 1818: data <= 'd0; 1819: data <= 'd0; 1820: data <= 'd0; 1821: data <= 'd0; 1822: data <= 'd0; 1823: data <= 'd0; 1824: data <= 'd0; 1825: data <= 'd0; 1826: data <= 'd0; 1827: data <= 'd0; 1828: data <= 'd0; 1829: data <= 'd0; 1830: data <= 'd0; 1831: data <= 'd0; 1832: data <= 'd0; 1833: data <= 'd0; 1834: data <= 'd2; 1835: data <= 'd9; 1836: data <= 'd9; 1837: data <= 'd2; 1838: data <= 'd1; 1839: data <= 'd3; 1840: data <= 'd3; 1841: data <= 'd1; 1842: data <= 'd1; 1843: data <= 'd3; 1844: data <= 'd1; 1845: data <= 'd1; 1846: data <= 'd2; 1847: data <= 'd0; 1848: data <= 'd0; 1849: data <= 'd0; 1850: data <= 'd0; 1851: data <= 'd0; 1852: data <= 'd0; 1853: data <= 'd0; 1854: data <= 'd0; 1855: data <= 'd0; 1856: data <= 'd0; 1857: data <= 'd0; 1858: data <= 'd0; 1859: data <= 'd0; 1860: data <= 'd0; 1861: data <= 'd0; 1862: data <= 'd0; 1863: data <= 'd0; 1864: data <= 'd0; 1865: data <= 'd0; 1866: data <= 'd2; 1867: data <= 'd9; 1868: data <= 'd9; 1869: data <= 'd2; 1870: data <= 'd2; 1871: data <= 'd2; 1872: data <= 'd5; 1873: data <= 'd5; 1874: data <= 'd5; 1875: data <= 'd2; 1876: data <= 'd2; 1877: data <= 'd2; 1878: data <= 'd2; 1879: data <= 'd0; 1880: data <= 'd0; 1881: data <= 'd0; 1882: data <= 'd0; 1883: data <= 'd0; 1884: data <= 'd0; 1885: data <= 'd0; 1886: data <= 'd0; 1887: data <= 'd0; 1888: data <= 'd0; 1889: data <= 'd0; 1890: data <= 'd0; 1891: data <= 'd0; 1892: data <= 'd0; 1893: data <= 'd0; 1894: data <= 'd0; 1895: data <= 'd0; 1896: data <= 'd0; 1897: data <= 'd0; 1898: data <= 'd0; 1899: data <= 'd2; 1900: data <= 'd2; 1901: data <= 'd1; 1902: data <= 'd3; 1903: data <= 'd3; 1904: data <= 'd3; 1905: data <= 'd1; 1906: data <= 'd3; 1907: data <= 'd3; 1908: data <= 'd3; 1909: data <= 'd5; 1910: data <= 'd2; 1911: data <= 'd0; 1912: data <= 'd0; 1913: data <= 'd0; 1914: data <= 'd0; 1915: data <= 'd0; 1916: data <= 'd0; 1917: data <= 'd0; 1918: data <= 'd0; 1919: data <= 'd0; 1920: data <= 'd0; 1921: data <= 'd0; 1922: data <= 'd0; 1923: data <= 'd0; 1924: data <= 'd0; 1925: data <= 'd0; 1926: data <= 'd0; 1927: data <= 'd0; 1928: data <= 'd0; 1929: data <= 'd0; 1930: data <= 'd0; 1931: data <= 'd2; 1932: data <= 'd4; 1933: data <= 'd7; 1934: data <= 'd7; 1935: data <= 'd2; 1936: data <= 'd2; 1937: data <= 'd2; 1938: data <= 'd2; 1939: data <= 'd5; 1940: data <= 'd5; 1941: data <= 'd4; 1942: data <= 'd2; 1943: data <= 'd0; 1944: data <= 'd0; 1945: data <= 'd0; 1946: data <= 'd0; 1947: data <= 'd0; 1948: data <= 'd0; 1949: data <= 'd0; 1950: data <= 'd0; 1951: data <= 'd0; 1952: data <= 'd0; 1953: data <= 'd0; 1954: data <= 'd0; 1955: data <= 'd0; 1956: data <= 'd0; 1957: data <= 'd0; 1958: data <= 'd0; 1959: data <= 'd0; 1960: data <= 'd0; 1961: data <= 'd0; 1962: data <= 'd0; 1963: data <= 'd2; 1964: data <= 'd4; 1965: data <= 'd7; 1966: data <= 'd2; 1967: data <= 'd0; 1968: data <= 'd0; 1969: data <= 'd0; 1970: data <= 'd0; 1971: data <= 'd2; 1972: data <= 'd4; 1973: data <= 'd4; 1974: data <= 'd2; 1975: data <= 'd0; 1976: data <= 'd0; 1977: data <= 'd0; 1978: data <= 'd0; 1979: data <= 'd0; 1980: data <= 'd0; 1981: data <= 'd0; 1982: data <= 'd0; 1983: data <= 'd0; 1984: data <= 'd0; 1985: data <= 'd0; 1986: data <= 'd0; 1987: data <= 'd0; 1988: data <= 'd0; 1989: data <= 'd0; 1990: data <= 'd0; 1991: data <= 'd0; 1992: data <= 'd0; 1993: data <= 'd0; 1994: data <= 'd0; 1995: data <= 'd2; 1996: data <= 'd2; 1997: data <= 'd2; 1998: data <= 'd0; 1999: data <= 'd0; 2000: data <= 'd0; 2001: data <= 'd0; 2002: data <= 'd0; 2003: data <= 'd0; 2004: data <= 'd2; 2005: data <= 'd2; 2006: data <= 'd2; 2007: data <= 'd0; 2008: data <= 'd0; 2009: data <= 'd0; 2010: data <= 'd0; 2011: data <= 'd0; 2012: data <= 'd0; 2013: data <= 'd0; 2014: data <= 'd0; 2015: data <= 'd0; 2016: data <= 'd0; 2017: data <= 'd0; 2018: data <= 'd0; 2019: data <= 'd0; 2020: data <= 'd0; 2021: data <= 'd0; 2022: data <= 'd0; 2023: data <= 'd0; 2024: data <= 'd0; 2025: data <= 'd0; 2026: data <= 'd0; 2027: data <= 'd0; 2028: data <= 'd0; 2029: data <= 'd0; 2030: data <= 'd0; 2031: data <= 'd0; 2032: data <= 'd0; 2033: data <= 'd0; 2034: data <= 'd0; 2035: data <= 'd0; 2036: data <= 'd0; 2037: data <= 'd0; 2038: data <= 'd0; 2039: data <= 'd0; 2040: data <= 'd0; 2041: data <= 'd0; 2042: data <= 'd0; 2043: data <= 'd0; 2044: data <= 'd0; 2045: data <= 'd0; 2046: data <= 'd0; 2047: data <= 'd0; 2048: data <= 'd0; 2049: data <= 'd0; 2050: data <= 'd0; 2051: data <= 'd0; 2052: data <= 'd0; 2053: data <= 'd0; 2054: data <= 'd0; 2055: data <= 'd0; 2056: data <= 'd0; 2057: data <= 'd0; 2058: data <= 'd0; 2059: data <= 'd0; 2060: data <= 'd0; 2061: data <= 'd0; 2062: data <= 'd0; 2063: data <= 'd0; 2064: data <= 'd0; 2065: data <= 'd0; 2066: data <= 'd0; 2067: data <= 'd0; 2068: data <= 'd0; 2069: data <= 'd0; 2070: data <= 'd0; 2071: data <= 'd0; 2072: data <= 'd0; 2073: data <= 'd0; 2074: data <= 'd0; 2075: data <= 'd0; 2076: data <= 'd0; 2077: data <= 'd0; 2078: data <= 'd0; 2079: data <= 'd0; 2080: data <= 'd0; 2081: data <= 'd0; 2082: data <= 'd0; 2083: data <= 'd0; 2084: data <= 'd0; 2085: data <= 'd0; 2086: data <= 'd0; 2087: data <= 'd0; 2088: data <= 'd0; 2089: data <= 'd0; 2090: data <= 'd0; 2091: data <= 'd0; 2092: data <= 'd0; 2093: data <= 'd0; 2094: data <= 'd0; 2095: data <= 'd0; 2096: data <= 'd0; 2097: data <= 'd0; 2098: data <= 'd0; 2099: data <= 'd0; 2100: data <= 'd0; 2101: data <= 'd0; 2102: data <= 'd0; 2103: data <= 'd0; 2104: data <= 'd0; 2105: data <= 'd0; 2106: data <= 'd0; 2107: data <= 'd0; 2108: data <= 'd0; 2109: data <= 'd0; 2110: data <= 'd0; 2111: data <= 'd0; 2112: data <= 'd0; 2113: data <= 'd0; 2114: data <= 'd0; 2115: data <= 'd0; 2116: data <= 'd0; 2117: data <= 'd0; 2118: data <= 'd0; 2119: data <= 'd0; 2120: data <= 'd0; 2121: data <= 'd0; 2122: data <= 'd0; 2123: data <= 'd0; 2124: data <= 'd0; 2125: data <= 'd0; 2126: data <= 'd0; 2127: data <= 'd0; 2128: data <= 'd0; 2129: data <= 'd0; 2130: data <= 'd0; 2131: data <= 'd0; 2132: data <= 'd0; 2133: data <= 'd0; 2134: data <= 'd0; 2135: data <= 'd0; 2136: data <= 'd0; 2137: data <= 'd0; 2138: data <= 'd0; 2139: data <= 'd0; 2140: data <= 'd0; 2141: data <= 'd0; 2142: data <= 'd0; 2143: data <= 'd0; 2144: data <= 'd0; 2145: data <= 'd0; 2146: data <= 'd0; 2147: data <= 'd0; 2148: data <= 'd0; 2149: data <= 'd0; 2150: data <= 'd0; 2151: data <= 'd0; 2152: data <= 'd0; 2153: data <= 'd0; 2154: data <= 'd0; 2155: data <= 'd0; 2156: data <= 'd0; 2157: data <= 'd0; 2158: data <= 'd0; 2159: data <= 'd0; 2160: data <= 'd0; 2161: data <= 'd0; 2162: data <= 'd0; 2163: data <= 'd0; 2164: data <= 'd0; 2165: data <= 'd0; 2166: data <= 'd0; 2167: data <= 'd0; 2168: data <= 'd0; 2169: data <= 'd0; 2170: data <= 'd0; 2171: data <= 'd0; 2172: data <= 'd0; 2173: data <= 'd0; 2174: data <= 'd0; 2175: data <= 'd0; 2176: data <= 'd0; 2177: data <= 'd0; 2178: data <= 'd0; 2179: data <= 'd0; 2180: data <= 'd0; 2181: data <= 'd0; 2182: data <= 'd0; 2183: data <= 'd0; 2184: data <= 'd0; 2185: data <= 'd0; 2186: data <= 'd0; 2187: data <= 'd0; 2188: data <= 'd0; 2189: data <= 'd0; 2190: data <= 'd0; 2191: data <= 'd0; 2192: data <= 'd0; 2193: data <= 'd0; 2194: data <= 'd0; 2195: data <= 'd0; 2196: data <= 'd0; 2197: data <= 'd0; 2198: data <= 'd0; 2199: data <= 'd0; 2200: data <= 'd0; 2201: data <= 'd0; 2202: data <= 'd0; 2203: data <= 'd0; 2204: data <= 'd0; 2205: data <= 'd0; 2206: data <= 'd0; 2207: data <= 'd0; 2208: data <= 'd0; 2209: data <= 'd0; 2210: data <= 'd0; 2211: data <= 'd0; 2212: data <= 'd0; 2213: data <= 'd0; 2214: data <= 'd0; 2215: data <= 'd0; 2216: data <= 'd0; 2217: data <= 'd0; 2218: data <= 'd0; 2219: data <= 'd0; 2220: data <= 'd0; 2221: data <= 'd0; 2222: data <= 'd0; 2223: data <= 'd0; 2224: data <= 'd0; 2225: data <= 'd0; 2226: data <= 'd0; 2227: data <= 'd0; 2228: data <= 'd0; 2229: data <= 'd0; 2230: data <= 'd0; 2231: data <= 'd0; 2232: data <= 'd0; 2233: data <= 'd0; 2234: data <= 'd0; 2235: data <= 'd0; 2236: data <= 'd0; 2237: data <= 'd0; 2238: data <= 'd0; 2239: data <= 'd0; 2240: data <= 'd0; 2241: data <= 'd0; 2242: data <= 'd0; 2243: data <= 'd0; 2244: data <= 'd0; 2245: data <= 'd0; 2246: data <= 'd0; 2247: data <= 'd0; 2248: data <= 'd0; 2249: data <= 'd0; 2250: data <= 'd0; 2251: data <= 'd0; 2252: data <= 'd0; 2253: data <= 'd0; 2254: data <= 'd0; 2255: data <= 'd0; 2256: data <= 'd0; 2257: data <= 'd0; 2258: data <= 'd0; 2259: data <= 'd0; 2260: data <= 'd0; 2261: data <= 'd0; 2262: data <= 'd0; 2263: data <= 'd0; 2264: data <= 'd0; 2265: data <= 'd0; 2266: data <= 'd0; 2267: data <= 'd0; 2268: data <= 'd0; 2269: data <= 'd0; 2270: data <= 'd0; 2271: data <= 'd0; 2272: data <= 'd0; 2273: data <= 'd0; 2274: data <= 'd0; 2275: data <= 'd0; 2276: data <= 'd0; 2277: data <= 'd0; 2278: data <= 'd0; 2279: data <= 'd0; 2280: data <= 'd0; 2281: data <= 'd0; 2282: data <= 'd0; 2283: data <= 'd0; 2284: data <= 'd0; 2285: data <= 'd0; 2286: data <= 'd0; 2287: data <= 'd0; 2288: data <= 'd0; 2289: data <= 'd0; 2290: data <= 'd0; 2291: data <= 'd0; 2292: data <= 'd0; 2293: data <= 'd0; 2294: data <= 'd0; 2295: data <= 'd0; 2296: data <= 'd0; 2297: data <= 'd0; 2298: data <= 'd0; 2299: data <= 'd0; 2300: data <= 'd0; 2301: data <= 'd0; 2302: data <= 'd0; 2303: data <= 'd0; 2304: data <= 'd0; 2305: data <= 'd0; 2306: data <= 'd0; 2307: data <= 'd0; 2308: data <= 'd0; 2309: data <= 'd0; 2310: data <= 'd0; 2311: data <= 'd0; 2312: data <= 'd0; 2313: data <= 'd0; 2314: data <= 'd0; 2315: data <= 'd0; 2316: data <= 'd0; 2317: data <= 'd0; 2318: data <= 'd0; 2319: data <= 'd0; 2320: data <= 'd0; 2321: data <= 'd0; 2322: data <= 'd0; 2323: data <= 'd0; 2324: data <= 'd0; 2325: data <= 'd0; 2326: data <= 'd0; 2327: data <= 'd0; 2328: data <= 'd0; 2329: data <= 'd0; 2330: data <= 'd0; 2331: data <= 'd0; 2332: data <= 'd0; 2333: data <= 'd0; 2334: data <= 'd0; 2335: data <= 'd0; 2336: data <= 'd0; 2337: data <= 'd0; 2338: data <= 'd0; 2339: data <= 'd0; 2340: data <= 'd0; 2341: data <= 'd0; 2342: data <= 'd0; 2343: data <= 'd0; 2344: data <= 'd0; 2345: data <= 'd0; 2346: data <= 'd0; 2347: data <= 'd0; 2348: data <= 'd0; 2349: data <= 'd2; 2350: data <= 'd2; 2351: data <= 'd2; 2352: data <= 'd2; 2353: data <= 'd2; 2354: data <= 'd2; 2355: data <= 'd0; 2356: data <= 'd0; 2357: data <= 'd0; 2358: data <= 'd0; 2359: data <= 'd0; 2360: data <= 'd0; 2361: data <= 'd0; 2362: data <= 'd0; 2363: data <= 'd0; 2364: data <= 'd0; 2365: data <= 'd0; 2366: data <= 'd0; 2367: data <= 'd0; 2368: data <= 'd0; 2369: data <= 'd0; 2370: data <= 'd0; 2371: data <= 'd0; 2372: data <= 'd0; 2373: data <= 'd0; 2374: data <= 'd0; 2375: data <= 'd0; 2376: data <= 'd0; 2377: data <= 'd0; 2378: data <= 'd0; 2379: data <= 'd2; 2380: data <= 'd2; 2381: data <= 'd6; 2382: data <= 'd6; 2383: data <= 'd6; 2384: data <= 'd6; 2385: data <= 'd6; 2386: data <= 'd6; 2387: data <= 'd2; 2388: data <= 'd2; 2389: data <= 'd0; 2390: data <= 'd0; 2391: data <= 'd0; 2392: data <= 'd0; 2393: data <= 'd0; 2394: data <= 'd0; 2395: data <= 'd0; 2396: data <= 'd0; 2397: data <= 'd0; 2398: data <= 'd0; 2399: data <= 'd0; 2400: data <= 'd0; 2401: data <= 'd0; 2402: data <= 'd0; 2403: data <= 'd0; 2404: data <= 'd0; 2405: data <= 'd0; 2406: data <= 'd0; 2407: data <= 'd0; 2408: data <= 'd0; 2409: data <= 'd0; 2410: data <= 'd2; 2411: data <= 'd1; 2412: data <= 'd3; 2413: data <= 'd6; 2414: data <= 'd6; 2415: data <= 'd6; 2416: data <= 'd6; 2417: data <= 'd6; 2418: data <= 'd6; 2419: data <= 'd6; 2420: data <= 'd3; 2421: data <= 'd2; 2422: data <= 'd0; 2423: data <= 'd0; 2424: data <= 'd0; 2425: data <= 'd0; 2426: data <= 'd0; 2427: data <= 'd0; 2428: data <= 'd0; 2429: data <= 'd0; 2430: data <= 'd0; 2431: data <= 'd0; 2432: data <= 'd0; 2433: data <= 'd0; 2434: data <= 'd0; 2435: data <= 'd0; 2436: data <= 'd0; 2437: data <= 'd0; 2438: data <= 'd0; 2439: data <= 'd0; 2440: data <= 'd0; 2441: data <= 'd2; 2442: data <= 'd1; 2443: data <= 'd1; 2444: data <= 'd1; 2445: data <= 'd3; 2446: data <= 'd6; 2447: data <= 'd6; 2448: data <= 'd6; 2449: data <= 'd6; 2450: data <= 'd6; 2451: data <= 'd3; 2452: data <= 'd1; 2453: data <= 'd1; 2454: data <= 'd2; 2455: data <= 'd0; 2456: data <= 'd0; 2457: data <= 'd0; 2458: data <= 'd0; 2459: data <= 'd0; 2460: data <= 'd0; 2461: data <= 'd0; 2462: data <= 'd0; 2463: data <= 'd0; 2464: data <= 'd0; 2465: data <= 'd0; 2466: data <= 'd0; 2467: data <= 'd0; 2468: data <= 'd0; 2469: data <= 'd0; 2470: data <= 'd0; 2471: data <= 'd0; 2472: data <= 'd0; 2473: data <= 'd2; 2474: data <= 'd1; 2475: data <= 'd1; 2476: data <= 'd5; 2477: data <= 'd5; 2478: data <= 'd5; 2479: data <= 'd1; 2480: data <= 'd1; 2481: data <= 'd1; 2482: data <= 'd1; 2483: data <= 'd1; 2484: data <= 'd5; 2485: data <= 'd5; 2486: data <= 'd2; 2487: data <= 'd0; 2488: data <= 'd0; 2489: data <= 'd0; 2490: data <= 'd0; 2491: data <= 'd0; 2492: data <= 'd0; 2493: data <= 'd0; 2494: data <= 'd0; 2495: data <= 'd0; 2496: data <= 'd0; 2497: data <= 'd0; 2498: data <= 'd0; 2499: data <= 'd0; 2500: data <= 'd0; 2501: data <= 'd0; 2502: data <= 'd0; 2503: data <= 'd0; 2504: data <= 'd2; 2505: data <= 'd1; 2506: data <= 'd5; 2507: data <= 'd5; 2508: data <= 'd3; 2509: data <= 'd6; 2510: data <= 'd6; 2511: data <= 'd6; 2512: data <= 'd6; 2513: data <= 'd6; 2514: data <= 'd6; 2515: data <= 'd6; 2516: data <= 'd6; 2517: data <= 'd3; 2518: data <= 'd5; 2519: data <= 'd2; 2520: data <= 'd0; 2521: data <= 'd0; 2522: data <= 'd0; 2523: data <= 'd0; 2524: data <= 'd0; 2525: data <= 'd0; 2526: data <= 'd0; 2527: data <= 'd0; 2528: data <= 'd0; 2529: data <= 'd0; 2530: data <= 'd0; 2531: data <= 'd0; 2532: data <= 'd0; 2533: data <= 'd0; 2534: data <= 'd0; 2535: data <= 'd0; 2536: data <= 'd2; 2537: data <= 'd5; 2538: data <= 'd3; 2539: data <= 'd6; 2540: data <= 'd3; 2541: data <= 'd1; 2542: data <= 'd1; 2543: data <= 'd1; 2544: data <= 'd1; 2545: data <= 'd1; 2546: data <= 'd1; 2547: data <= 'd1; 2548: data <= 'd1; 2549: data <= 'd1; 2550: data <= 'd3; 2551: data <= 'd2; 2552: data <= 'd0; 2553: data <= 'd0; 2554: data <= 'd0; 2555: data <= 'd0; 2556: data <= 'd0; 2557: data <= 'd0; 2558: data <= 'd0; 2559: data <= 'd0; 2560: data <= 'd0; 2561: data <= 'd0; 2562: data <= 'd0; 2563: data <= 'd0; 2564: data <= 'd0; 2565: data <= 'd0; 2566: data <= 'd0; 2567: data <= 'd0; 2568: data <= 'd2; 2569: data <= 'd5; 2570: data <= 'd3; 2571: data <= 'd1; 2572: data <= 'd1; 2573: data <= 'd1; 2574: data <= 'd5; 2575: data <= 'd5; 2576: data <= 'd5; 2577: data <= 'd5; 2578: data <= 'd5; 2579: data <= 'd5; 2580: data <= 'd5; 2581: data <= 'd1; 2582: data <= 'd1; 2583: data <= 'd2; 2584: data <= 'd0; 2585: data <= 'd0; 2586: data <= 'd0; 2587: data <= 'd0; 2588: data <= 'd0; 2589: data <= 'd0; 2590: data <= 'd0; 2591: data <= 'd0; 2592: data <= 'd0; 2593: data <= 'd0; 2594: data <= 'd0; 2595: data <= 'd0; 2596: data <= 'd0; 2597: data <= 'd0; 2598: data <= 'd0; 2599: data <= 'd0; 2600: data <= 'd2; 2601: data <= 'd6; 2602: data <= 'd1; 2603: data <= 'd5; 2604: data <= 'd2; 2605: data <= 'd2; 2606: data <= 'd2; 2607: data <= 'd2; 2608: data <= 'd2; 2609: data <= 'd2; 2610: data <= 'd2; 2611: data <= 'd2; 2612: data <= 'd2; 2613: data <= 'd2; 2614: data <= 'd5; 2615: data <= 'd2; 2616: data <= 'd0; 2617: data <= 'd0; 2618: data <= 'd0; 2619: data <= 'd0; 2620: data <= 'd0; 2621: data <= 'd0; 2622: data <= 'd0; 2623: data <= 'd0; 2624: data <= 'd0; 2625: data <= 'd0; 2626: data <= 'd0; 2627: data <= 'd0; 2628: data <= 'd0; 2629: data <= 'd0; 2630: data <= 'd2; 2631: data <= 'd2; 2632: data <= 'd2; 2633: data <= 'd1; 2634: data <= 'd5; 2635: data <= 'd2; 2636: data <= 'd8; 2637: data <= 'd8; 2638: data <= 'd8; 2639: data <= 'd8; 2640: data <= 'd8; 2641: data <= 'd9; 2642: data <= 'd9; 2643: data <= 'd8; 2644: data <= 'd8; 2645: data <= 'd8; 2646: data <= 'd2; 2647: data <= 'd2; 2648: data <= 'd0; 2649: data <= 'd0; 2650: data <= 'd0; 2651: data <= 'd0; 2652: data <= 'd0; 2653: data <= 'd0; 2654: data <= 'd0; 2655: data <= 'd0; 2656: data <= 'd0; 2657: data <= 'd0; 2658: data <= 'd0; 2659: data <= 'd0; 2660: data <= 'd0; 2661: data <= 'd0; 2662: data <= 'd2; 2663: data <= 'd1; 2664: data <= 'd2; 2665: data <= 'd1; 2666: data <= 'd2; 2667: data <= 'd8; 2668: data <= 'd8; 2669: data <= 'd9; 2670: data <= 'd9; 2671: data <= 'd2; 2672: data <= 'd9; 2673: data <= 'd11; 2674: data <= 'd11; 2675: data <= 'd10; 2676: data <= 'd2; 2677: data <= 'd9; 2678: data <= 'd2; 2679: data <= 'd2; 2680: data <= 'd0; 2681: data <= 'd0; 2682: data <= 'd0; 2683: data <= 'd0; 2684: data <= 'd0; 2685: data <= 'd0; 2686: data <= 'd0; 2687: data <= 'd0; 2688: data <= 'd0; 2689: data <= 'd0; 2690: data <= 'd0; 2691: data <= 'd0; 2692: data <= 'd0; 2693: data <= 'd0; 2694: data <= 'd2; 2695: data <= 'd5; 2696: data <= 'd1; 2697: data <= 'd2; 2698: data <= 'd9; 2699: data <= 'd10; 2700: data <= 'd9; 2701: data <= 'd9; 2702: data <= 'd10; 2703: data <= 'd11; 2704: data <= 'd10; 2705: data <= 'd11; 2706: data <= 'd11; 2707: data <= 'd10; 2708: data <= 'd11; 2709: data <= 'd10; 2710: data <= 'd9; 2711: data <= 'd2; 2712: data <= 'd0; 2713: data <= 'd0; 2714: data <= 'd0; 2715: data <= 'd0; 2716: data <= 'd0; 2717: data <= 'd0; 2718: data <= 'd0; 2719: data <= 'd0; 2720: data <= 'd0; 2721: data <= 'd0; 2722: data <= 'd0; 2723: data <= 'd0; 2724: data <= 'd0; 2725: data <= 'd0; 2726: data <= 'd0; 2727: data <= 'd2; 2728: data <= 'd5; 2729: data <= 'd5; 2730: data <= 'd2; 2731: data <= 'd8; 2732: data <= 'd9; 2733: data <= 'd9; 2734: data <= 'd10; 2735: data <= 'd10; 2736: data <= 'd10; 2737: data <= 'd8; 2738: data <= 'd8; 2739: data <= 'd10; 2740: data <= 'd10; 2741: data <= 'd9; 2742: data <= 'd2; 2743: data <= 'd0; 2744: data <= 'd0; 2745: data <= 'd0; 2746: data <= 'd0; 2747: data <= 'd0; 2748: data <= 'd0; 2749: data <= 'd0; 2750: data <= 'd0; 2751: data <= 'd0; 2752: data <= 'd0; 2753: data <= 'd0; 2754: data <= 'd0; 2755: data <= 'd0; 2756: data <= 'd0; 2757: data <= 'd0; 2758: data <= 'd0; 2759: data <= 'd0; 2760: data <= 'd2; 2761: data <= 'd2; 2762: data <= 'd2; 2763: data <= 'd8; 2764: data <= 'd8; 2765: data <= 'd9; 2766: data <= 'd9; 2767: data <= 'd10; 2768: data <= 'd10; 2769: data <= 'd9; 2770: data <= 'd9; 2771: data <= 'd10; 2772: data <= 'd10; 2773: data <= 'd9; 2774: data <= 'd2; 2775: data <= 'd0; 2776: data <= 'd0; 2777: data <= 'd0; 2778: data <= 'd0; 2779: data <= 'd0; 2780: data <= 'd0; 2781: data <= 'd0; 2782: data <= 'd0; 2783: data <= 'd0; 2784: data <= 'd0; 2785: data <= 'd0; 2786: data <= 'd0; 2787: data <= 'd0; 2788: data <= 'd0; 2789: data <= 'd0; 2790: data <= 'd0; 2791: data <= 'd0; 2792: data <= 'd0; 2793: data <= 'd0; 2794: data <= 'd2; 2795: data <= 'd2; 2796: data <= 'd5; 2797: data <= 'd5; 2798: data <= 'd8; 2799: data <= 'd9; 2800: data <= 'd9; 2801: data <= 'd9; 2802: data <= 'd9; 2803: data <= 'd9; 2804: data <= 'd9; 2805: data <= 'd5; 2806: data <= 'd2; 2807: data <= 'd0; 2808: data <= 'd0; 2809: data <= 'd0; 2810: data <= 'd0; 2811: data <= 'd0; 2812: data <= 'd0; 2813: data <= 'd0; 2814: data <= 'd0; 2815: data <= 'd0; 2816: data <= 'd0; 2817: data <= 'd0; 2818: data <= 'd0; 2819: data <= 'd0; 2820: data <= 'd0; 2821: data <= 'd0; 2822: data <= 'd0; 2823: data <= 'd0; 2824: data <= 'd0; 2825: data <= 'd2; 2826: data <= 'd7; 2827: data <= 'd1; 2828: data <= 'd1; 2829: data <= 'd1; 2830: data <= 'd3; 2831: data <= 'd3; 2832: data <= 'd3; 2833: data <= 'd5; 2834: data <= 'd5; 2835: data <= 'd3; 2836: data <= 'd3; 2837: data <= 'd1; 2838: data <= 'd2; 2839: data <= 'd0; 2840: data <= 'd0; 2841: data <= 'd0; 2842: data <= 'd0; 2843: data <= 'd0; 2844: data <= 'd0; 2845: data <= 'd0; 2846: data <= 'd0; 2847: data <= 'd0; 2848: data <= 'd0; 2849: data <= 'd0; 2850: data <= 'd0; 2851: data <= 'd0; 2852: data <= 'd0; 2853: data <= 'd0; 2854: data <= 'd0; 2855: data <= 'd0; 2856: data <= 'd0; 2857: data <= 'd2; 2858: data <= 'd7; 2859: data <= 'd7; 2860: data <= 'd1; 2861: data <= 'd1; 2862: data <= 'd3; 2863: data <= 'd3; 2864: data <= 'd3; 2865: data <= 'd1; 2866: data <= 'd1; 2867: data <= 'd3; 2868: data <= 'd3; 2869: data <= 'd1; 2870: data <= 'd2; 2871: data <= 'd0; 2872: data <= 'd0; 2873: data <= 'd0; 2874: data <= 'd0; 2875: data <= 'd0; 2876: data <= 'd0; 2877: data <= 'd0; 2878: data <= 'd0; 2879: data <= 'd0; 2880: data <= 'd0; 2881: data <= 'd0; 2882: data <= 'd0; 2883: data <= 'd0; 2884: data <= 'd0; 2885: data <= 'd0; 2886: data <= 'd0; 2887: data <= 'd0; 2888: data <= 'd2; 2889: data <= 'd9; 2890: data <= 'd9; 2891: data <= 'd7; 2892: data <= 'd1; 2893: data <= 'd1; 2894: data <= 'd1; 2895: data <= 'd3; 2896: data <= 'd3; 2897: data <= 'd1; 2898: data <= 'd1; 2899: data <= 'd3; 2900: data <= 'd1; 2901: data <= 'd1; 2902: data <= 'd8; 2903: data <= 'd2; 2904: data <= 'd0; 2905: data <= 'd0; 2906: data <= 'd0; 2907: data <= 'd0; 2908: data <= 'd0; 2909: data <= 'd0; 2910: data <= 'd0; 2911: data <= 'd0; 2912: data <= 'd0; 2913: data <= 'd0; 2914: data <= 'd0; 2915: data <= 'd0; 2916: data <= 'd0; 2917: data <= 'd0; 2918: data <= 'd0; 2919: data <= 'd0; 2920: data <= 'd2; 2921: data <= 'd9; 2922: data <= 'd9; 2923: data <= 'd2; 2924: data <= 'd2; 2925: data <= 'd2; 2926: data <= 'd2; 2927: data <= 'd2; 2928: data <= 'd5; 2929: data <= 'd5; 2930: data <= 'd5; 2931: data <= 'd2; 2932: data <= 'd2; 2933: data <= 'd2; 2934: data <= 'd8; 2935: data <= 'd2; 2936: data <= 'd0; 2937: data <= 'd0; 2938: data <= 'd0; 2939: data <= 'd0; 2940: data <= 'd0; 2941: data <= 'd0; 2942: data <= 'd0; 2943: data <= 'd0; 2944: data <= 'd0; 2945: data <= 'd0; 2946: data <= 'd0; 2947: data <= 'd0; 2948: data <= 'd0; 2949: data <= 'd0; 2950: data <= 'd0; 2951: data <= 'd0; 2952: data <= 'd0; 2953: data <= 'd2; 2954: data <= 'd2; 2955: data <= 'd2; 2956: data <= 'd1; 2957: data <= 'd1; 2958: data <= 'd3; 2959: data <= 'd3; 2960: data <= 'd3; 2961: data <= 'd1; 2962: data <= 'd3; 2963: data <= 'd3; 2964: data <= 'd3; 2965: data <= 'd2; 2966: data <= 'd2; 2967: data <= 'd0; 2968: data <= 'd0; 2969: data <= 'd0; 2970: data <= 'd0; 2971: data <= 'd0; 2972: data <= 'd0; 2973: data <= 'd0; 2974: data <= 'd0; 2975: data <= 'd0; 2976: data <= 'd0; 2977: data <= 'd0; 2978: data <= 'd0; 2979: data <= 'd0; 2980: data <= 'd0; 2981: data <= 'd0; 2982: data <= 'd0; 2983: data <= 'd0; 2984: data <= 'd0; 2985: data <= 'd0; 2986: data <= 'd0; 2987: data <= 'd2; 2988: data <= 'd4; 2989: data <= 'd7; 2990: data <= 'd7; 2991: data <= 'd2; 2992: data <= 'd2; 2993: data <= 'd2; 2994: data <= 'd5; 2995: data <= 'd5; 2996: data <= 'd4; 2997: data <= 'd2; 2998: data <= 'd0; 2999: data <= 'd0; 3000: data <= 'd0; 3001: data <= 'd0; 3002: data <= 'd0; 3003: data <= 'd0; 3004: data <= 'd0; 3005: data <= 'd0; 3006: data <= 'd0; 3007: data <= 'd0; 3008: data <= 'd0; 3009: data <= 'd0; 3010: data <= 'd0; 3011: data <= 'd0; 3012: data <= 'd0; 3013: data <= 'd0; 3014: data <= 'd0; 3015: data <= 'd0; 3016: data <= 'd0; 3017: data <= 'd0; 3018: data <= 'd0; 3019: data <= 'd2; 3020: data <= 'd4; 3021: data <= 'd7; 3022: data <= 'd2; 3023: data <= 'd0; 3024: data <= 'd0; 3025: data <= 'd0; 3026: data <= 'd2; 3027: data <= 'd4; 3028: data <= 'd4; 3029: data <= 'd2; 3030: data <= 'd0; 3031: data <= 'd0; 3032: data <= 'd0; 3033: data <= 'd0; 3034: data <= 'd0; 3035: data <= 'd0; 3036: data <= 'd0; 3037: data <= 'd0; 3038: data <= 'd0; 3039: data <= 'd0; 3040: data <= 'd0; 3041: data <= 'd0; 3042: data <= 'd0; 3043: data <= 'd0; 3044: data <= 'd0; 3045: data <= 'd0; 3046: data <= 'd0; 3047: data <= 'd0; 3048: data <= 'd0; 3049: data <= 'd0; 3050: data <= 'd0; 3051: data <= 'd2; 3052: data <= 'd2; 3053: data <= 'd2; 3054: data <= 'd0; 3055: data <= 'd0; 3056: data <= 'd0; 3057: data <= 'd0; 3058: data <= 'd2; 3059: data <= 'd2; 3060: data <= 'd2; 3061: data <= 'd0; 3062: data <= 'd0; 3063: data <= 'd0; 3064: data <= 'd0; 3065: data <= 'd0; 3066: data <= 'd0; 3067: data <= 'd0; 3068: data <= 'd0; 3069: data <= 'd0; 3070: data <= 'd0; 3071: data <= 'd0; 3072: data <= 'd0; 3073: data <= 'd0; 3074: data <= 'd0; 3075: data <= 'd0; 3076: data <= 'd0; 3077: data <= 'd0; 3078: data <= 'd0; 3079: data <= 'd0; 3080: data <= 'd0; 3081: data <= 'd0; 3082: data <= 'd0; 3083: data <= 'd0; 3084: data <= 'd0; 3085: data <= 'd0; 3086: data <= 'd0; 3087: data <= 'd0; 3088: data <= 'd0; 3089: data <= 'd0; 3090: data <= 'd0; 3091: data <= 'd0; 3092: data <= 'd0; 3093: data <= 'd0; 3094: data <= 'd0; 3095: data <= 'd0; 3096: data <= 'd0; 3097: data <= 'd0; 3098: data <= 'd0; 3099: data <= 'd0; 3100: data <= 'd0; 3101: data <= 'd0; 3102: data <= 'd0; 3103: data <= 'd0; 3104: data <= 'd0; 3105: data <= 'd0; 3106: data <= 'd0; 3107: data <= 'd0; 3108: data <= 'd0; 3109: data <= 'd0; 3110: data <= 'd0; 3111: data <= 'd0; 3112: data <= 'd0; 3113: data <= 'd0; 3114: data <= 'd0; 3115: data <= 'd0; 3116: data <= 'd0; 3117: data <= 'd0; 3118: data <= 'd0; 3119: data <= 'd0; 3120: data <= 'd0; 3121: data <= 'd0; 3122: data <= 'd0; 3123: data <= 'd0; 3124: data <= 'd0; 3125: data <= 'd0; 3126: data <= 'd0; 3127: data <= 'd0; 3128: data <= 'd0; 3129: data <= 'd0; 3130: data <= 'd0; 3131: data <= 'd0; 3132: data <= 'd0; 3133: data <= 'd0; 3134: data <= 'd0; 3135: data <= 'd0; 3136: data <= 'd0; 3137: data <= 'd0; 3138: data <= 'd0; 3139: data <= 'd0; 3140: data <= 'd0; 3141: data <= 'd0; 3142: data <= 'd0; 3143: data <= 'd0; 3144: data <= 'd0; 3145: data <= 'd0; 3146: data <= 'd0; 3147: data <= 'd0; 3148: data <= 'd0; 3149: data <= 'd0; 3150: data <= 'd0; 3151: data <= 'd0; 3152: data <= 'd0; 3153: data <= 'd0; 3154: data <= 'd0; 3155: data <= 'd0; 3156: data <= 'd0; 3157: data <= 'd0; 3158: data <= 'd0; 3159: data <= 'd0; 3160: data <= 'd0; 3161: data <= 'd0; 3162: data <= 'd0; 3163: data <= 'd0; 3164: data <= 'd0; 3165: data <= 'd0; 3166: data <= 'd0; 3167: data <= 'd0; 3168: data <= 'd0; 3169: data <= 'd0; 3170: data <= 'd0; 3171: data <= 'd0; 3172: data <= 'd0; 3173: data <= 'd0; 3174: data <= 'd0; 3175: data <= 'd0; 3176: data <= 'd0; 3177: data <= 'd0; 3178: data <= 'd0; 3179: data <= 'd0; 3180: data <= 'd0; 3181: data <= 'd0; 3182: data <= 'd0; 3183: data <= 'd0; 3184: data <= 'd0; 3185: data <= 'd0; 3186: data <= 'd0; 3187: data <= 'd0; 3188: data <= 'd0; 3189: data <= 'd0; 3190: data <= 'd0; 3191: data <= 'd0; 3192: data <= 'd0; 3193: data <= 'd0; 3194: data <= 'd0; 3195: data <= 'd0; 3196: data <= 'd0; 3197: data <= 'd0; 3198: data <= 'd0; 3199: data <= 'd0; 3200: data <= 'd0; 3201: data <= 'd0; 3202: data <= 'd0; 3203: data <= 'd0; 3204: data <= 'd0; 3205: data <= 'd0; 3206: data <= 'd0; 3207: data <= 'd0; 3208: data <= 'd0; 3209: data <= 'd0; 3210: data <= 'd0; 3211: data <= 'd0; 3212: data <= 'd0; 3213: data <= 'd0; 3214: data <= 'd0; 3215: data <= 'd0; 3216: data <= 'd0; 3217: data <= 'd0; 3218: data <= 'd0; 3219: data <= 'd0; 3220: data <= 'd0; 3221: data <= 'd0; 3222: data <= 'd0; 3223: data <= 'd0; 3224: data <= 'd0; 3225: data <= 'd0; 3226: data <= 'd0; 3227: data <= 'd0; 3228: data <= 'd0; 3229: data <= 'd0; 3230: data <= 'd0; 3231: data <= 'd0; 3232: data <= 'd0; 3233: data <= 'd0; 3234: data <= 'd0; 3235: data <= 'd0; 3236: data <= 'd0; 3237: data <= 'd0; 3238: data <= 'd0; 3239: data <= 'd0; 3240: data <= 'd0; 3241: data <= 'd0; 3242: data <= 'd0; 3243: data <= 'd0; 3244: data <= 'd0; 3245: data <= 'd0; 3246: data <= 'd0; 3247: data <= 'd0; 3248: data <= 'd0; 3249: data <= 'd0; 3250: data <= 'd0; 3251: data <= 'd0; 3252: data <= 'd0; 3253: data <= 'd0; 3254: data <= 'd0; 3255: data <= 'd0; 3256: data <= 'd0; 3257: data <= 'd0; 3258: data <= 'd0; 3259: data <= 'd0; 3260: data <= 'd0; 3261: data <= 'd0; 3262: data <= 'd0; 3263: data <= 'd0; 3264: data <= 'd0; 3265: data <= 'd0; 3266: data <= 'd0; 3267: data <= 'd0; 3268: data <= 'd0; 3269: data <= 'd0; 3270: data <= 'd0; 3271: data <= 'd0; 3272: data <= 'd0; 3273: data <= 'd0; 3274: data <= 'd0; 3275: data <= 'd0; 3276: data <= 'd0; 3277: data <= 'd0; 3278: data <= 'd0; 3279: data <= 'd0; 3280: data <= 'd0; 3281: data <= 'd0; 3282: data <= 'd0; 3283: data <= 'd0; 3284: data <= 'd0; 3285: data <= 'd0; 3286: data <= 'd0; 3287: data <= 'd0; 3288: data <= 'd0; 3289: data <= 'd0; 3290: data <= 'd0; 3291: data <= 'd0; 3292: data <= 'd0; 3293: data <= 'd0; 3294: data <= 'd0; 3295: data <= 'd0; 3296: data <= 'd0; 3297: data <= 'd0; 3298: data <= 'd0; 3299: data <= 'd0; 3300: data <= 'd0; 3301: data <= 'd0; 3302: data <= 'd0; 3303: data <= 'd0; 3304: data <= 'd0; 3305: data <= 'd0; 3306: data <= 'd0; 3307: data <= 'd0; 3308: data <= 'd0; 3309: data <= 'd0; 3310: data <= 'd0; 3311: data <= 'd0; 3312: data <= 'd0; 3313: data <= 'd0; 3314: data <= 'd0; 3315: data <= 'd0; 3316: data <= 'd0; 3317: data <= 'd0; 3318: data <= 'd0; 3319: data <= 'd0; 3320: data <= 'd0; 3321: data <= 'd0; 3322: data <= 'd0; 3323: data <= 'd0; 3324: data <= 'd0; 3325: data <= 'd0; 3326: data <= 'd0; 3327: data <= 'd0; 3328: data <= 'd0; 3329: data <= 'd0; 3330: data <= 'd0; 3331: data <= 'd0; 3332: data <= 'd0; 3333: data <= 'd0; 3334: data <= 'd0; 3335: data <= 'd0; 3336: data <= 'd0; 3337: data <= 'd0; 3338: data <= 'd0; 3339: data <= 'd0; 3340: data <= 'd0; 3341: data <= 'd2; 3342: data <= 'd2; 3343: data <= 'd2; 3344: data <= 'd2; 3345: data <= 'd2; 3346: data <= 'd2; 3347: data <= 'd0; 3348: data <= 'd0; 3349: data <= 'd0; 3350: data <= 'd0; 3351: data <= 'd0; 3352: data <= 'd0; 3353: data <= 'd0; 3354: data <= 'd0; 3355: data <= 'd0; 3356: data <= 'd0; 3357: data <= 'd0; 3358: data <= 'd0; 3359: data <= 'd0; 3360: data <= 'd0; 3361: data <= 'd0; 3362: data <= 'd0; 3363: data <= 'd0; 3364: data <= 'd0; 3365: data <= 'd0; 3366: data <= 'd0; 3367: data <= 'd0; 3368: data <= 'd0; 3369: data <= 'd0; 3370: data <= 'd0; 3371: data <= 'd2; 3372: data <= 'd2; 3373: data <= 'd6; 3374: data <= 'd6; 3375: data <= 'd6; 3376: data <= 'd6; 3377: data <= 'd6; 3378: data <= 'd6; 3379: data <= 'd2; 3380: data <= 'd2; 3381: data <= 'd0; 3382: data <= 'd0; 3383: data <= 'd0; 3384: data <= 'd0; 3385: data <= 'd0; 3386: data <= 'd0; 3387: data <= 'd0; 3388: data <= 'd0; 3389: data <= 'd0; 3390: data <= 'd0; 3391: data <= 'd0; 3392: data <= 'd0; 3393: data <= 'd0; 3394: data <= 'd0; 3395: data <= 'd0; 3396: data <= 'd0; 3397: data <= 'd0; 3398: data <= 'd0; 3399: data <= 'd0; 3400: data <= 'd0; 3401: data <= 'd0; 3402: data <= 'd2; 3403: data <= 'd1; 3404: data <= 'd3; 3405: data <= 'd6; 3406: data <= 'd6; 3407: data <= 'd6; 3408: data <= 'd6; 3409: data <= 'd6; 3410: data <= 'd6; 3411: data <= 'd6; 3412: data <= 'd3; 3413: data <= 'd2; 3414: data <= 'd0; 3415: data <= 'd0; 3416: data <= 'd0; 3417: data <= 'd0; 3418: data <= 'd0; 3419: data <= 'd0; 3420: data <= 'd0; 3421: data <= 'd0; 3422: data <= 'd0; 3423: data <= 'd0; 3424: data <= 'd0; 3425: data <= 'd0; 3426: data <= 'd0; 3427: data <= 'd0; 3428: data <= 'd0; 3429: data <= 'd0; 3430: data <= 'd0; 3431: data <= 'd0; 3432: data <= 'd0; 3433: data <= 'd2; 3434: data <= 'd1; 3435: data <= 'd1; 3436: data <= 'd1; 3437: data <= 'd3; 3438: data <= 'd6; 3439: data <= 'd6; 3440: data <= 'd6; 3441: data <= 'd6; 3442: data <= 'd6; 3443: data <= 'd3; 3444: data <= 'd1; 3445: data <= 'd1; 3446: data <= 'd2; 3447: data <= 'd0; 3448: data <= 'd0; 3449: data <= 'd0; 3450: data <= 'd0; 3451: data <= 'd0; 3452: data <= 'd0; 3453: data <= 'd0; 3454: data <= 'd0; 3455: data <= 'd0; 3456: data <= 'd0; 3457: data <= 'd0; 3458: data <= 'd0; 3459: data <= 'd0; 3460: data <= 'd0; 3461: data <= 'd0; 3462: data <= 'd0; 3463: data <= 'd0; 3464: data <= 'd0; 3465: data <= 'd2; 3466: data <= 'd1; 3467: data <= 'd1; 3468: data <= 'd5; 3469: data <= 'd5; 3470: data <= 'd5; 3471: data <= 'd1; 3472: data <= 'd1; 3473: data <= 'd1; 3474: data <= 'd1; 3475: data <= 'd1; 3476: data <= 'd5; 3477: data <= 'd5; 3478: data <= 'd2; 3479: data <= 'd0; 3480: data <= 'd0; 3481: data <= 'd0; 3482: data <= 'd0; 3483: data <= 'd0; 3484: data <= 'd0; 3485: data <= 'd0; 3486: data <= 'd0; 3487: data <= 'd0; 3488: data <= 'd0; 3489: data <= 'd0; 3490: data <= 'd0; 3491: data <= 'd0; 3492: data <= 'd0; 3493: data <= 'd0; 3494: data <= 'd0; 3495: data <= 'd0; 3496: data <= 'd2; 3497: data <= 'd1; 3498: data <= 'd5; 3499: data <= 'd5; 3500: data <= 'd3; 3501: data <= 'd6; 3502: data <= 'd6; 3503: data <= 'd6; 3504: data <= 'd6; 3505: data <= 'd6; 3506: data <= 'd6; 3507: data <= 'd6; 3508: data <= 'd6; 3509: data <= 'd3; 3510: data <= 'd5; 3511: data <= 'd2; 3512: data <= 'd0; 3513: data <= 'd0; 3514: data <= 'd0; 3515: data <= 'd0; 3516: data <= 'd0; 3517: data <= 'd0; 3518: data <= 'd0; 3519: data <= 'd0; 3520: data <= 'd0; 3521: data <= 'd0; 3522: data <= 'd0; 3523: data <= 'd0; 3524: data <= 'd0; 3525: data <= 'd0; 3526: data <= 'd0; 3527: data <= 'd0; 3528: data <= 'd2; 3529: data <= 'd5; 3530: data <= 'd3; 3531: data <= 'd6; 3532: data <= 'd3; 3533: data <= 'd1; 3534: data <= 'd1; 3535: data <= 'd1; 3536: data <= 'd1; 3537: data <= 'd1; 3538: data <= 'd1; 3539: data <= 'd1; 3540: data <= 'd1; 3541: data <= 'd1; 3542: data <= 'd3; 3543: data <= 'd2; 3544: data <= 'd0; 3545: data <= 'd0; 3546: data <= 'd0; 3547: data <= 'd0; 3548: data <= 'd0; 3549: data <= 'd0; 3550: data <= 'd0; 3551: data <= 'd0; 3552: data <= 'd0; 3553: data <= 'd0; 3554: data <= 'd0; 3555: data <= 'd0; 3556: data <= 'd0; 3557: data <= 'd0; 3558: data <= 'd0; 3559: data <= 'd0; 3560: data <= 'd2; 3561: data <= 'd5; 3562: data <= 'd3; 3563: data <= 'd1; 3564: data <= 'd1; 3565: data <= 'd1; 3566: data <= 'd5; 3567: data <= 'd5; 3568: data <= 'd5; 3569: data <= 'd5; 3570: data <= 'd5; 3571: data <= 'd5; 3572: data <= 'd5; 3573: data <= 'd1; 3574: data <= 'd1; 3575: data <= 'd2; 3576: data <= 'd0; 3577: data <= 'd0; 3578: data <= 'd0; 3579: data <= 'd0; 3580: data <= 'd0; 3581: data <= 'd0; 3582: data <= 'd0; 3583: data <= 'd0; 3584: data <= 'd0; 3585: data <= 'd0; 3586: data <= 'd0; 3587: data <= 'd0; 3588: data <= 'd0; 3589: data <= 'd0; 3590: data <= 'd0; 3591: data <= 'd0; 3592: data <= 'd2; 3593: data <= 'd6; 3594: data <= 'd1; 3595: data <= 'd5; 3596: data <= 'd2; 3597: data <= 'd2; 3598: data <= 'd2; 3599: data <= 'd2; 3600: data <= 'd2; 3601: data <= 'd2; 3602: data <= 'd2; 3603: data <= 'd2; 3604: data <= 'd2; 3605: data <= 'd2; 3606: data <= 'd5; 3607: data <= 'd2; 3608: data <= 'd0; 3609: data <= 'd0; 3610: data <= 'd0; 3611: data <= 'd0; 3612: data <= 'd0; 3613: data <= 'd0; 3614: data <= 'd0; 3615: data <= 'd0; 3616: data <= 'd0; 3617: data <= 'd0; 3618: data <= 'd0; 3619: data <= 'd0; 3620: data <= 'd0; 3621: data <= 'd0; 3622: data <= 'd2; 3623: data <= 'd2; 3624: data <= 'd5; 3625: data <= 'd6; 3626: data <= 'd5; 3627: data <= 'd2; 3628: data <= 'd8; 3629: data <= 'd8; 3630: data <= 'd8; 3631: data <= 'd8; 3632: data <= 'd8; 3633: data <= 'd9; 3634: data <= 'd9; 3635: data <= 'd8; 3636: data <= 'd8; 3637: data <= 'd8; 3638: data <= 'd2; 3639: data <= 'd2; 3640: data <= 'd0; 3641: data <= 'd0; 3642: data <= 'd0; 3643: data <= 'd0; 3644: data <= 'd0; 3645: data <= 'd0; 3646: data <= 'd0; 3647: data <= 'd0; 3648: data <= 'd0; 3649: data <= 'd0; 3650: data <= 'd0; 3651: data <= 'd0; 3652: data <= 'd0; 3653: data <= 'd0; 3654: data <= 'd2; 3655: data <= 'd3; 3656: data <= 'd6; 3657: data <= 'd3; 3658: data <= 'd2; 3659: data <= 'd8; 3660: data <= 'd8; 3661: data <= 'd9; 3662: data <= 'd9; 3663: data <= 'd10; 3664: data <= 'd2; 3665: data <= 'd9; 3666: data <= 'd11; 3667: data <= 'd10; 3668: data <= 'd2; 3669: data <= 'd9; 3670: data <= 'd2; 3671: data <= 'd2; 3672: data <= 'd0; 3673: data <= 'd0; 3674: data <= 'd0; 3675: data <= 'd0; 3676: data <= 'd0; 3677: data <= 'd0; 3678: data <= 'd0; 3679: data <= 'd0; 3680: data <= 'd0; 3681: data <= 'd0; 3682: data <= 'd0; 3683: data <= 'd0; 3684: data <= 'd0; 3685: data <= 'd0; 3686: data <= 'd2; 3687: data <= 'd1; 3688: data <= 'd3; 3689: data <= 'd1; 3690: data <= 'd2; 3691: data <= 'd10; 3692: data <= 'd10; 3693: data <= 'd9; 3694: data <= 'd10; 3695: data <= 'd10; 3696: data <= 'd11; 3697: data <= 'd10; 3698: data <= 'd11; 3699: data <= 'd11; 3700: data <= 'd10; 3701: data <= 'd10; 3702: data <= 'd2; 3703: data <= 'd0; 3704: data <= 'd0; 3705: data <= 'd0; 3706: data <= 'd0; 3707: data <= 'd0; 3708: data <= 'd0; 3709: data <= 'd0; 3710: data <= 'd0; 3711: data <= 'd0; 3712: data <= 'd0; 3713: data <= 'd0; 3714: data <= 'd0; 3715: data <= 'd0; 3716: data <= 'd0; 3717: data <= 'd0; 3718: data <= 'd0; 3719: data <= 'd2; 3720: data <= 'd1; 3721: data <= 'd5; 3722: data <= 'd2; 3723: data <= 'd8; 3724: data <= 'd9; 3725: data <= 'd9; 3726: data <= 'd10; 3727: data <= 'd10; 3728: data <= 'd10; 3729: data <= 'd10; 3730: data <= 'd8; 3731: data <= 'd8; 3732: data <= 'd10; 3733: data <= 'd9; 3734: data <= 'd2; 3735: data <= 'd0; 3736: data <= 'd0; 3737: data <= 'd0; 3738: data <= 'd0; 3739: data <= 'd0; 3740: data <= 'd0; 3741: data <= 'd0; 3742: data <= 'd0; 3743: data <= 'd0; 3744: data <= 'd0; 3745: data <= 'd0; 3746: data <= 'd0; 3747: data <= 'd0; 3748: data <= 'd0; 3749: data <= 'd0; 3750: data <= 'd0; 3751: data <= 'd0; 3752: data <= 'd2; 3753: data <= 'd2; 3754: data <= 'd2; 3755: data <= 'd8; 3756: data <= 'd8; 3757: data <= 'd9; 3758: data <= 'd9; 3759: data <= 'd10; 3760: data <= 'd10; 3761: data <= 'd10; 3762: data <= 'd9; 3763: data <= 'd9; 3764: data <= 'd10; 3765: data <= 'd9; 3766: data <= 'd2; 3767: data <= 'd0; 3768: data <= 'd0; 3769: data <= 'd0; 3770: data <= 'd0; 3771: data <= 'd0; 3772: data <= 'd0; 3773: data <= 'd0; 3774: data <= 'd0; 3775: data <= 'd0; 3776: data <= 'd0; 3777: data <= 'd0; 3778: data <= 'd0; 3779: data <= 'd0; 3780: data <= 'd0; 3781: data <= 'd0; 3782: data <= 'd0; 3783: data <= 'd0; 3784: data <= 'd0; 3785: data <= 'd0; 3786: data <= 'd0; 3787: data <= 'd2; 3788: data <= 'd5; 3789: data <= 'd5; 3790: data <= 'd8; 3791: data <= 'd9; 3792: data <= 'd9; 3793: data <= 'd9; 3794: data <= 'd9; 3795: data <= 'd9; 3796: data <= 'd9; 3797: data <= 'd2; 3798: data <= 'd0; 3799: data <= 'd0; 3800: data <= 'd0; 3801: data <= 'd0; 3802: data <= 'd0; 3803: data <= 'd0; 3804: data <= 'd0; 3805: data <= 'd0; 3806: data <= 'd0; 3807: data <= 'd0; 3808: data <= 'd0; 3809: data <= 'd0; 3810: data <= 'd0; 3811: data <= 'd0; 3812: data <= 'd0; 3813: data <= 'd0; 3814: data <= 'd0; 3815: data <= 'd0; 3816: data <= 'd0; 3817: data <= 'd0; 3818: data <= 'd2; 3819: data <= 'd7; 3820: data <= 'd1; 3821: data <= 'd1; 3822: data <= 'd1; 3823: data <= 'd3; 3824: data <= 'd3; 3825: data <= 'd3; 3826: data <= 'd5; 3827: data <= 'd5; 3828: data <= 'd3; 3829: data <= 'd1; 3830: data <= 'd2; 3831: data <= 'd0; 3832: data <= 'd0; 3833: data <= 'd0; 3834: data <= 'd0; 3835: data <= 'd0; 3836: data <= 'd0; 3837: data <= 'd0; 3838: data <= 'd0; 3839: data <= 'd0; 3840: data <= 'd0; 3841: data <= 'd0; 3842: data <= 'd0; 3843: data <= 'd0; 3844: data <= 'd0; 3845: data <= 'd0; 3846: data <= 'd0; 3847: data <= 'd0; 3848: data <= 'd0; 3849: data <= 'd2; 3850: data <= 'd7; 3851: data <= 'd7; 3852: data <= 'd7; 3853: data <= 'd1; 3854: data <= 'd1; 3855: data <= 'd3; 3856: data <= 'd3; 3857: data <= 'd3; 3858: data <= 'd1; 3859: data <= 'd1; 3860: data <= 'd3; 3861: data <= 'd1; 3862: data <= 'd2; 3863: data <= 'd2; 3864: data <= 'd0; 3865: data <= 'd0; 3866: data <= 'd0; 3867: data <= 'd0; 3868: data <= 'd0; 3869: data <= 'd0; 3870: data <= 'd0; 3871: data <= 'd0; 3872: data <= 'd0; 3873: data <= 'd0; 3874: data <= 'd0; 3875: data <= 'd0; 3876: data <= 'd0; 3877: data <= 'd0; 3878: data <= 'd0; 3879: data <= 'd0; 3880: data <= 'd2; 3881: data <= 'd8; 3882: data <= 'd10; 3883: data <= 'd10; 3884: data <= 'd5; 3885: data <= 'd1; 3886: data <= 'd1; 3887: data <= 'd1; 3888: data <= 'd3; 3889: data <= 'd3; 3890: data <= 'd1; 3891: data <= 'd1; 3892: data <= 'd1; 3893: data <= 'd1; 3894: data <= 'd8; 3895: data <= 'd9; 3896: data <= 'd2; 3897: data <= 'd0; 3898: data <= 'd0; 3899: data <= 'd0; 3900: data <= 'd0; 3901: data <= 'd0; 3902: data <= 'd0; 3903: data <= 'd0; 3904: data <= 'd0; 3905: data <= 'd0; 3906: data <= 'd0; 3907: data <= 'd0; 3908: data <= 'd0; 3909: data <= 'd0; 3910: data <= 'd0; 3911: data <= 'd0; 3912: data <= 'd2; 3913: data <= 'd9; 3914: data <= 'd10; 3915: data <= 'd9; 3916: data <= 'd2; 3917: data <= 'd2; 3918: data <= 'd2; 3919: data <= 'd2; 3920: data <= 'd2; 3921: data <= 'd5; 3922: data <= 'd5; 3923: data <= 'd5; 3924: data <= 'd2; 3925: data <= 'd2; 3926: data <= 'd8; 3927: data <= 'd9; 3928: data <= 'd2; 3929: data <= 'd0; 3930: data <= 'd0; 3931: data <= 'd0; 3932: data <= 'd0; 3933: data <= 'd0; 3934: data <= 'd0; 3935: data <= 'd0; 3936: data <= 'd0; 3937: data <= 'd0; 3938: data <= 'd0; 3939: data <= 'd0; 3940: data <= 'd0; 3941: data <= 'd0; 3942: data <= 'd0; 3943: data <= 'd0; 3944: data <= 'd0; 3945: data <= 'd2; 3946: data <= 'd2; 3947: data <= 'd2; 3948: data <= 'd2; 3949: data <= 'd1; 3950: data <= 'd1; 3951: data <= 'd3; 3952: data <= 'd3; 3953: data <= 'd3; 3954: data <= 'd1; 3955: data <= 'd3; 3956: data <= 'd3; 3957: data <= 'd2; 3958: data <= 'd2; 3959: data <= 'd2; 3960: data <= 'd0; 3961: data <= 'd0; 3962: data <= 'd0; 3963: data <= 'd0; 3964: data <= 'd0; 3965: data <= 'd0; 3966: data <= 'd0; 3967: data <= 'd0; 3968: data <= 'd0; 3969: data <= 'd0; 3970: data <= 'd0; 3971: data <= 'd0; 3972: data <= 'd0; 3973: data <= 'd0; 3974: data <= 'd0; 3975: data <= 'd0; 3976: data <= 'd0; 3977: data <= 'd0; 3978: data <= 'd0; 3979: data <= 'd2; 3980: data <= 'd4; 3981: data <= 'd7; 3982: data <= 'd7; 3983: data <= 'd2; 3984: data <= 'd2; 3985: data <= 'd2; 3986: data <= 'd5; 3987: data <= 'd5; 3988: data <= 'd4; 3989: data <= 'd2; 3990: data <= 'd0; 3991: data <= 'd0; 3992: data <= 'd0; 3993: data <= 'd0; 3994: data <= 'd0; 3995: data <= 'd0; 3996: data <= 'd0; 3997: data <= 'd0; 3998: data <= 'd0; 3999: data <= 'd0; 4000: data <= 'd0; 4001: data <= 'd0; 4002: data <= 'd0; 4003: data <= 'd0; 4004: data <= 'd0; 4005: data <= 'd0; 4006: data <= 'd0; 4007: data <= 'd0; 4008: data <= 'd0; 4009: data <= 'd0; 4010: data <= 'd0; 4011: data <= 'd0; 4012: data <= 'd2; 4013: data <= 'd4; 4014: data <= 'd7; 4015: data <= 'd2; 4016: data <= 'd0; 4017: data <= 'd2; 4018: data <= 'd4; 4019: data <= 'd4; 4020: data <= 'd2; 4021: data <= 'd0; 4022: data <= 'd0; 4023: data <= 'd0; 4024: data <= 'd0; 4025: data <= 'd0; 4026: data <= 'd0; 4027: data <= 'd0; 4028: data <= 'd0; 4029: data <= 'd0; 4030: data <= 'd0; 4031: data <= 'd0; 4032: data <= 'd0; 4033: data <= 'd0; 4034: data <= 'd0; 4035: data <= 'd0; 4036: data <= 'd0; 4037: data <= 'd0; 4038: data <= 'd0; 4039: data <= 'd0; 4040: data <= 'd0; 4041: data <= 'd0; 4042: data <= 'd0; 4043: data <= 'd0; 4044: data <= 'd0; 4045: data <= 'd2; 4046: data <= 'd2; 4047: data <= 'd2; 4048: data <= 'd0; 4049: data <= 'd2; 4050: data <= 'd2; 4051: data <= 'd2; 4052: data <= 'd0; 4053: data <= 'd0; 4054: data <= 'd0; 4055: data <= 'd0; 4056: data <= 'd0; 4057: data <= 'd0; 4058: data <= 'd0; 4059: data <= 'd0; 4060: data <= 'd0; 4061: data <= 'd0; 4062: data <= 'd0; 4063: data <= 'd0; 4064: data <= 'd0; 4065: data <= 'd0; 4066: data <= 'd0; 4067: data <= 'd0; 4068: data <= 'd0; 4069: data <= 'd0; 4070: data <= 'd0; 4071: data <= 'd0; 4072: data <= 'd0; 4073: data <= 'd0; 4074: data <= 'd0; 4075: data <= 'd0; 4076: data <= 'd0; 4077: data <= 'd0; 4078: data <= 'd0; 4079: data <= 'd0; 4080: data <= 'd0; 4081: data <= 'd0; 4082: data <= 'd0; 4083: data <= 'd0; 4084: data <= 'd0; 4085: data <= 'd0; 4086: data <= 'd0; 4087: data <= 'd0; 4088: data <= 'd0; 4089: data <= 'd0; 4090: data <= 'd0; 4091: data <= 'd0; 4092: data <= 'd0; 4093: data <= 'd0; 4094: data <= 'd0; 4095: data <= 'd0; 4096: data <= 'd0; 4097: data <= 'd0; 4098: data <= 'd0; 4099: data <= 'd0; 4100: data <= 'd0; 4101: data <= 'd0; 4102: data <= 'd0; 4103: data <= 'd0; 4104: data <= 'd0; 4105: data <= 'd0; 4106: data <= 'd0; 4107: data <= 'd0; 4108: data <= 'd0; 4109: data <= 'd0; 4110: data <= 'd0; 4111: data <= 'd0; 4112: data <= 'd0; 4113: data <= 'd0; 4114: data <= 'd0; 4115: data <= 'd0; 4116: data <= 'd0; 4117: data <= 'd0; 4118: data <= 'd0; 4119: data <= 'd0; 4120: data <= 'd0; 4121: data <= 'd0; 4122: data <= 'd0; 4123: data <= 'd0; 4124: data <= 'd0; 4125: data <= 'd0; 4126: data <= 'd0; 4127: data <= 'd0; 4128: data <= 'd0; 4129: data <= 'd0; 4130: data <= 'd0; 4131: data <= 'd0; 4132: data <= 'd0; 4133: data <= 'd0; 4134: data <= 'd0; 4135: data <= 'd0; 4136: data <= 'd0; 4137: data <= 'd0; 4138: data <= 'd0; 4139: data <= 'd0; 4140: data <= 'd0; 4141: data <= 'd0; 4142: data <= 'd0; 4143: data <= 'd0; 4144: data <= 'd0; 4145: data <= 'd0; 4146: data <= 'd0; 4147: data <= 'd0; 4148: data <= 'd0; 4149: data <= 'd0; 4150: data <= 'd0; 4151: data <= 'd0; 4152: data <= 'd0; 4153: data <= 'd0; 4154: data <= 'd0; 4155: data <= 'd0; 4156: data <= 'd0; 4157: data <= 'd0; 4158: data <= 'd0; 4159: data <= 'd0; 4160: data <= 'd0; 4161: data <= 'd0; 4162: data <= 'd0; 4163: data <= 'd0; 4164: data <= 'd0; 4165: data <= 'd0; 4166: data <= 'd0; 4167: data <= 'd0; 4168: data <= 'd0; 4169: data <= 'd0; 4170: data <= 'd0; 4171: data <= 'd0; 4172: data <= 'd0; 4173: data <= 'd0; 4174: data <= 'd0; 4175: data <= 'd0; 4176: data <= 'd0; 4177: data <= 'd0; 4178: data <= 'd0; 4179: data <= 'd0; 4180: data <= 'd0; 4181: data <= 'd0; 4182: data <= 'd0; 4183: data <= 'd0; 4184: data <= 'd0; 4185: data <= 'd0; 4186: data <= 'd0; 4187: data <= 'd0; 4188: data <= 'd0; 4189: data <= 'd0; 4190: data <= 'd0; 4191: data <= 'd0; 4192: data <= 'd0; 4193: data <= 'd0; 4194: data <= 'd0; 4195: data <= 'd0; 4196: data <= 'd0; 4197: data <= 'd0; 4198: data <= 'd0; 4199: data <= 'd0; 4200: data <= 'd0; 4201: data <= 'd0; 4202: data <= 'd0; 4203: data <= 'd0; 4204: data <= 'd0; 4205: data <= 'd0; 4206: data <= 'd0; 4207: data <= 'd0; 4208: data <= 'd0; 4209: data <= 'd0; 4210: data <= 'd0; 4211: data <= 'd0; 4212: data <= 'd0; 4213: data <= 'd0; 4214: data <= 'd0; 4215: data <= 'd0; 4216: data <= 'd0; 4217: data <= 'd0; 4218: data <= 'd0; 4219: data <= 'd0; 4220: data <= 'd0; 4221: data <= 'd0; 4222: data <= 'd0; 4223: data <= 'd0; 4224: data <= 'd0; 4225: data <= 'd0; 4226: data <= 'd0; 4227: data <= 'd0; 4228: data <= 'd0; 4229: data <= 'd0; 4230: data <= 'd0; 4231: data <= 'd0; 4232: data <= 'd0; 4233: data <= 'd0; 4234: data <= 'd0; 4235: data <= 'd0; 4236: data <= 'd0; 4237: data <= 'd0; 4238: data <= 'd0; 4239: data <= 'd0; 4240: data <= 'd0; 4241: data <= 'd0; 4242: data <= 'd0; 4243: data <= 'd0; 4244: data <= 'd0; 4245: data <= 'd0; 4246: data <= 'd0; 4247: data <= 'd0; 4248: data <= 'd0; 4249: data <= 'd0; 4250: data <= 'd0; 4251: data <= 'd0; 4252: data <= 'd0; 4253: data <= 'd0; 4254: data <= 'd0; 4255: data <= 'd0; 4256: data <= 'd0; 4257: data <= 'd0; 4258: data <= 'd0; 4259: data <= 'd0; 4260: data <= 'd0; 4261: data <= 'd0; 4262: data <= 'd0; 4263: data <= 'd0; 4264: data <= 'd0; 4265: data <= 'd0; 4266: data <= 'd0; 4267: data <= 'd0; 4268: data <= 'd0; 4269: data <= 'd0; 4270: data <= 'd0; 4271: data <= 'd0; 4272: data <= 'd0; 4273: data <= 'd0; 4274: data <= 'd0; 4275: data <= 'd0; 4276: data <= 'd0; 4277: data <= 'd0; 4278: data <= 'd0; 4279: data <= 'd0; 4280: data <= 'd0; 4281: data <= 'd0; 4282: data <= 'd0; 4283: data <= 'd0; 4284: data <= 'd0; 4285: data <= 'd0; 4286: data <= 'd0; 4287: data <= 'd0; 4288: data <= 'd0; 4289: data <= 'd0; 4290: data <= 'd0; 4291: data <= 'd0; 4292: data <= 'd0; 4293: data <= 'd0; 4294: data <= 'd0; 4295: data <= 'd0; 4296: data <= 'd0; 4297: data <= 'd0; 4298: data <= 'd0; 4299: data <= 'd0; 4300: data <= 'd0; 4301: data <= 'd0; 4302: data <= 'd0; 4303: data <= 'd0; 4304: data <= 'd0; 4305: data <= 'd0; 4306: data <= 'd0; 4307: data <= 'd0; 4308: data <= 'd0; 4309: data <= 'd0; 4310: data <= 'd0; 4311: data <= 'd0; 4312: data <= 'd0; 4313: data <= 'd0; 4314: data <= 'd0; 4315: data <= 'd0; 4316: data <= 'd0; 4317: data <= 'd0; 4318: data <= 'd0; 4319: data <= 'd0; 4320: data <= 'd0; 4321: data <= 'd0; 4322: data <= 'd0; 4323: data <= 'd0; 4324: data <= 'd0; 4325: data <= 'd0; 4326: data <= 'd0; 4327: data <= 'd0; 4328: data <= 'd0; 4329: data <= 'd0; 4330: data <= 'd0; 4331: data <= 'd0; 4332: data <= 'd0; 4333: data <= 'd0; 4334: data <= 'd0; 4335: data <= 'd0; 4336: data <= 'd0; 4337: data <= 'd0; 4338: data <= 'd0; 4339: data <= 'd0; 4340: data <= 'd0; 4341: data <= 'd0; 4342: data <= 'd0; 4343: data <= 'd0; 4344: data <= 'd0; 4345: data <= 'd0; 4346: data <= 'd0; 4347: data <= 'd0; 4348: data <= 'd0; 4349: data <= 'd0; 4350: data <= 'd0; 4351: data <= 'd0; 4352: data <= 'd0; 4353: data <= 'd0; 4354: data <= 'd0; 4355: data <= 'd0; 4356: data <= 'd0; 4357: data <= 'd0; 4358: data <= 'd0; 4359: data <= 'd0; 4360: data <= 'd0; 4361: data <= 'd0; 4362: data <= 'd0; 4363: data <= 'd0; 4364: data <= 'd0; 4365: data <= 'd0; 4366: data <= 'd0; 4367: data <= 'd0; 4368: data <= 'd0; 4369: data <= 'd0; 4370: data <= 'd0; 4371: data <= 'd0; 4372: data <= 'd0; 4373: data <= 'd0; 4374: data <= 'd0; 4375: data <= 'd0; 4376: data <= 'd0; 4377: data <= 'd0; 4378: data <= 'd0; 4379: data <= 'd0; 4380: data <= 'd0; 4381: data <= 'd0; 4382: data <= 'd0; 4383: data <= 'd0; 4384: data <= 'd0; 4385: data <= 'd0; 4386: data <= 'd0; 4387: data <= 'd0; 4388: data <= 'd0; 4389: data <= 'd0; 4390: data <= 'd0; 4391: data <= 'd0; 4392: data <= 'd0; 4393: data <= 'd0; 4394: data <= 'd0; 4395: data <= 'd0; 4396: data <= 'd0; 4397: data <= 'd0; 4398: data <= 'd0; 4399: data <= 'd0; 4400: data <= 'd0; 4401: data <= 'd0; 4402: data <= 'd0; 4403: data <= 'd0; 4404: data <= 'd0; 4405: data <= 'd0; 4406: data <= 'd0; 4407: data <= 'd0; 4408: data <= 'd0; 4409: data <= 'd0; 4410: data <= 'd0; 4411: data <= 'd0; 4412: data <= 'd0; 4413: data <= 'd0; 4414: data <= 'd0; 4415: data <= 'd0; 4416: data <= 'd0; 4417: data <= 'd0; 4418: data <= 'd0; 4419: data <= 'd0; 4420: data <= 'd0; 4421: data <= 'd0; 4422: data <= 'd0; 4423: data <= 'd0; 4424: data <= 'd0; 4425: data <= 'd0; 4426: data <= 'd0; 4427: data <= 'd0; 4428: data <= 'd0; 4429: data <= 'd0; 4430: data <= 'd2; 4431: data <= 'd2; 4432: data <= 'd2; 4433: data <= 'd2; 4434: data <= 'd2; 4435: data <= 'd2; 4436: data <= 'd0; 4437: data <= 'd0; 4438: data <= 'd0; 4439: data <= 'd0; 4440: data <= 'd0; 4441: data <= 'd0; 4442: data <= 'd0; 4443: data <= 'd0; 4444: data <= 'd0; 4445: data <= 'd0; 4446: data <= 'd0; 4447: data <= 'd0; 4448: data <= 'd0; 4449: data <= 'd0; 4450: data <= 'd0; 4451: data <= 'd0; 4452: data <= 'd0; 4453: data <= 'd0; 4454: data <= 'd0; 4455: data <= 'd0; 4456: data <= 'd0; 4457: data <= 'd0; 4458: data <= 'd0; 4459: data <= 'd0; 4460: data <= 'd2; 4461: data <= 'd2; 4462: data <= 'd6; 4463: data <= 'd6; 4464: data <= 'd6; 4465: data <= 'd6; 4466: data <= 'd6; 4467: data <= 'd6; 4468: data <= 'd2; 4469: data <= 'd2; 4470: data <= 'd0; 4471: data <= 'd0; 4472: data <= 'd0; 4473: data <= 'd0; 4474: data <= 'd0; 4475: data <= 'd0; 4476: data <= 'd0; 4477: data <= 'd0; 4478: data <= 'd0; 4479: data <= 'd0; 4480: data <= 'd0; 4481: data <= 'd0; 4482: data <= 'd0; 4483: data <= 'd0; 4484: data <= 'd0; 4485: data <= 'd0; 4486: data <= 'd0; 4487: data <= 'd0; 4488: data <= 'd0; 4489: data <= 'd0; 4490: data <= 'd0; 4491: data <= 'd2; 4492: data <= 'd1; 4493: data <= 'd3; 4494: data <= 'd6; 4495: data <= 'd6; 4496: data <= 'd6; 4497: data <= 'd6; 4498: data <= 'd6; 4499: data <= 'd6; 4500: data <= 'd6; 4501: data <= 'd3; 4502: data <= 'd2; 4503: data <= 'd0; 4504: data <= 'd0; 4505: data <= 'd0; 4506: data <= 'd0; 4507: data <= 'd0; 4508: data <= 'd0; 4509: data <= 'd0; 4510: data <= 'd0; 4511: data <= 'd0; 4512: data <= 'd0; 4513: data <= 'd0; 4514: data <= 'd0; 4515: data <= 'd0; 4516: data <= 'd0; 4517: data <= 'd0; 4518: data <= 'd0; 4519: data <= 'd0; 4520: data <= 'd0; 4521: data <= 'd0; 4522: data <= 'd2; 4523: data <= 'd1; 4524: data <= 'd1; 4525: data <= 'd1; 4526: data <= 'd3; 4527: data <= 'd6; 4528: data <= 'd6; 4529: data <= 'd6; 4530: data <= 'd6; 4531: data <= 'd6; 4532: data <= 'd3; 4533: data <= 'd1; 4534: data <= 'd1; 4535: data <= 'd2; 4536: data <= 'd0; 4537: data <= 'd0; 4538: data <= 'd0; 4539: data <= 'd0; 4540: data <= 'd0; 4541: data <= 'd0; 4542: data <= 'd0; 4543: data <= 'd0; 4544: data <= 'd0; 4545: data <= 'd0; 4546: data <= 'd0; 4547: data <= 'd0; 4548: data <= 'd0; 4549: data <= 'd0; 4550: data <= 'd0; 4551: data <= 'd0; 4552: data <= 'd0; 4553: data <= 'd0; 4554: data <= 'd2; 4555: data <= 'd1; 4556: data <= 'd1; 4557: data <= 'd5; 4558: data <= 'd5; 4559: data <= 'd5; 4560: data <= 'd1; 4561: data <= 'd1; 4562: data <= 'd1; 4563: data <= 'd1; 4564: data <= 'd1; 4565: data <= 'd5; 4566: data <= 'd5; 4567: data <= 'd2; 4568: data <= 'd0; 4569: data <= 'd0; 4570: data <= 'd0; 4571: data <= 'd0; 4572: data <= 'd0; 4573: data <= 'd0; 4574: data <= 'd0; 4575: data <= 'd0; 4576: data <= 'd0; 4577: data <= 'd0; 4578: data <= 'd0; 4579: data <= 'd0; 4580: data <= 'd0; 4581: data <= 'd0; 4582: data <= 'd0; 4583: data <= 'd0; 4584: data <= 'd0; 4585: data <= 'd2; 4586: data <= 'd1; 4587: data <= 'd5; 4588: data <= 'd5; 4589: data <= 'd3; 4590: data <= 'd6; 4591: data <= 'd6; 4592: data <= 'd6; 4593: data <= 'd6; 4594: data <= 'd6; 4595: data <= 'd6; 4596: data <= 'd6; 4597: data <= 'd6; 4598: data <= 'd3; 4599: data <= 'd5; 4600: data <= 'd2; 4601: data <= 'd0; 4602: data <= 'd0; 4603: data <= 'd0; 4604: data <= 'd0; 4605: data <= 'd0; 4606: data <= 'd0; 4607: data <= 'd0; 4608: data <= 'd0; 4609: data <= 'd0; 4610: data <= 'd0; 4611: data <= 'd0; 4612: data <= 'd0; 4613: data <= 'd0; 4614: data <= 'd0; 4615: data <= 'd0; 4616: data <= 'd0; 4617: data <= 'd2; 4618: data <= 'd5; 4619: data <= 'd3; 4620: data <= 'd6; 4621: data <= 'd3; 4622: data <= 'd1; 4623: data <= 'd1; 4624: data <= 'd1; 4625: data <= 'd1; 4626: data <= 'd1; 4627: data <= 'd1; 4628: data <= 'd1; 4629: data <= 'd1; 4630: data <= 'd1; 4631: data <= 'd3; 4632: data <= 'd2; 4633: data <= 'd0; 4634: data <= 'd0; 4635: data <= 'd0; 4636: data <= 'd0; 4637: data <= 'd0; 4638: data <= 'd0; 4639: data <= 'd0; 4640: data <= 'd0; 4641: data <= 'd0; 4642: data <= 'd0; 4643: data <= 'd0; 4644: data <= 'd0; 4645: data <= 'd0; 4646: data <= 'd0; 4647: data <= 'd0; 4648: data <= 'd0; 4649: data <= 'd2; 4650: data <= 'd5; 4651: data <= 'd3; 4652: data <= 'd1; 4653: data <= 'd1; 4654: data <= 'd1; 4655: data <= 'd5; 4656: data <= 'd5; 4657: data <= 'd5; 4658: data <= 'd5; 4659: data <= 'd5; 4660: data <= 'd5; 4661: data <= 'd5; 4662: data <= 'd1; 4663: data <= 'd1; 4664: data <= 'd2; 4665: data <= 'd0; 4666: data <= 'd0; 4667: data <= 'd0; 4668: data <= 'd0; 4669: data <= 'd0; 4670: data <= 'd0; 4671: data <= 'd0; 4672: data <= 'd0; 4673: data <= 'd0; 4674: data <= 'd0; 4675: data <= 'd0; 4676: data <= 'd0; 4677: data <= 'd0; 4678: data <= 'd0; 4679: data <= 'd0; 4680: data <= 'd0; 4681: data <= 'd2; 4682: data <= 'd6; 4683: data <= 'd1; 4684: data <= 'd5; 4685: data <= 'd2; 4686: data <= 'd2; 4687: data <= 'd2; 4688: data <= 'd2; 4689: data <= 'd2; 4690: data <= 'd2; 4691: data <= 'd2; 4692: data <= 'd2; 4693: data <= 'd2; 4694: data <= 'd2; 4695: data <= 'd5; 4696: data <= 'd2; 4697: data <= 'd0; 4698: data <= 'd0; 4699: data <= 'd0; 4700: data <= 'd0; 4701: data <= 'd0; 4702: data <= 'd0; 4703: data <= 'd0; 4704: data <= 'd0; 4705: data <= 'd0; 4706: data <= 'd0; 4707: data <= 'd0; 4708: data <= 'd0; 4709: data <= 'd0; 4710: data <= 'd0; 4711: data <= 'd2; 4712: data <= 'd2; 4713: data <= 'd2; 4714: data <= 'd1; 4715: data <= 'd5; 4716: data <= 'd2; 4717: data <= 'd8; 4718: data <= 'd8; 4719: data <= 'd8; 4720: data <= 'd8; 4721: data <= 'd8; 4722: data <= 'd9; 4723: data <= 'd9; 4724: data <= 'd8; 4725: data <= 'd8; 4726: data <= 'd8; 4727: data <= 'd2; 4728: data <= 'd2; 4729: data <= 'd0; 4730: data <= 'd0; 4731: data <= 'd0; 4732: data <= 'd0; 4733: data <= 'd0; 4734: data <= 'd0; 4735: data <= 'd0; 4736: data <= 'd0; 4737: data <= 'd0; 4738: data <= 'd0; 4739: data <= 'd0; 4740: data <= 'd0; 4741: data <= 'd0; 4742: data <= 'd0; 4743: data <= 'd2; 4744: data <= 'd1; 4745: data <= 'd2; 4746: data <= 'd1; 4747: data <= 'd2; 4748: data <= 'd8; 4749: data <= 'd8; 4750: data <= 'd9; 4751: data <= 'd9; 4752: data <= 'd2; 4753: data <= 'd9; 4754: data <= 'd11; 4755: data <= 'd11; 4756: data <= 'd10; 4757: data <= 'd2; 4758: data <= 'd9; 4759: data <= 'd2; 4760: data <= 'd2; 4761: data <= 'd0; 4762: data <= 'd0; 4763: data <= 'd0; 4764: data <= 'd0; 4765: data <= 'd0; 4766: data <= 'd0; 4767: data <= 'd0; 4768: data <= 'd0; 4769: data <= 'd0; 4770: data <= 'd0; 4771: data <= 'd0; 4772: data <= 'd0; 4773: data <= 'd0; 4774: data <= 'd0; 4775: data <= 'd2; 4776: data <= 'd5; 4777: data <= 'd1; 4778: data <= 'd2; 4779: data <= 'd9; 4780: data <= 'd10; 4781: data <= 'd9; 4782: data <= 'd9; 4783: data <= 'd10; 4784: data <= 'd11; 4785: data <= 'd10; 4786: data <= 'd11; 4787: data <= 'd11; 4788: data <= 'd10; 4789: data <= 'd11; 4790: data <= 'd10; 4791: data <= 'd9; 4792: data <= 'd2; 4793: data <= 'd0; 4794: data <= 'd0; 4795: data <= 'd0; 4796: data <= 'd0; 4797: data <= 'd0; 4798: data <= 'd0; 4799: data <= 'd0; 4800: data <= 'd0; 4801: data <= 'd0; 4802: data <= 'd0; 4803: data <= 'd0; 4804: data <= 'd0; 4805: data <= 'd0; 4806: data <= 'd0; 4807: data <= 'd0; 4808: data <= 'd2; 4809: data <= 'd5; 4810: data <= 'd5; 4811: data <= 'd2; 4812: data <= 'd8; 4813: data <= 'd9; 4814: data <= 'd9; 4815: data <= 'd10; 4816: data <= 'd10; 4817: data <= 'd10; 4818: data <= 'd8; 4819: data <= 'd8; 4820: data <= 'd10; 4821: data <= 'd10; 4822: data <= 'd9; 4823: data <= 'd2; 4824: data <= 'd0; 4825: data <= 'd0; 4826: data <= 'd0; 4827: data <= 'd0; 4828: data <= 'd0; 4829: data <= 'd0; 4830: data <= 'd0; 4831: data <= 'd0; 4832: data <= 'd0; 4833: data <= 'd0; 4834: data <= 'd0; 4835: data <= 'd0; 4836: data <= 'd0; 4837: data <= 'd0; 4838: data <= 'd0; 4839: data <= 'd0; 4840: data <= 'd0; 4841: data <= 'd2; 4842: data <= 'd2; 4843: data <= 'd2; 4844: data <= 'd8; 4845: data <= 'd8; 4846: data <= 'd9; 4847: data <= 'd9; 4848: data <= 'd10; 4849: data <= 'd10; 4850: data <= 'd9; 4851: data <= 'd9; 4852: data <= 'd10; 4853: data <= 'd10; 4854: data <= 'd9; 4855: data <= 'd2; 4856: data <= 'd0; 4857: data <= 'd0; 4858: data <= 'd0; 4859: data <= 'd0; 4860: data <= 'd0; 4861: data <= 'd0; 4862: data <= 'd0; 4863: data <= 'd0; 4864: data <= 'd0; 4865: data <= 'd0; 4866: data <= 'd0; 4867: data <= 'd0; 4868: data <= 'd0; 4869: data <= 'd0; 4870: data <= 'd0; 4871: data <= 'd0; 4872: data <= 'd0; 4873: data <= 'd0; 4874: data <= 'd0; 4875: data <= 'd2; 4876: data <= 'd2; 4877: data <= 'd5; 4878: data <= 'd5; 4879: data <= 'd8; 4880: data <= 'd9; 4881: data <= 'd9; 4882: data <= 'd9; 4883: data <= 'd9; 4884: data <= 'd9; 4885: data <= 'd9; 4886: data <= 'd5; 4887: data <= 'd2; 4888: data <= 'd0; 4889: data <= 'd0; 4890: data <= 'd0; 4891: data <= 'd0; 4892: data <= 'd0; 4893: data <= 'd0; 4894: data <= 'd0; 4895: data <= 'd0; 4896: data <= 'd0; 4897: data <= 'd0; 4898: data <= 'd0; 4899: data <= 'd0; 4900: data <= 'd0; 4901: data <= 'd0; 4902: data <= 'd0; 4903: data <= 'd0; 4904: data <= 'd0; 4905: data <= 'd0; 4906: data <= 'd2; 4907: data <= 'd7; 4908: data <= 'd1; 4909: data <= 'd1; 4910: data <= 'd1; 4911: data <= 'd3; 4912: data <= 'd3; 4913: data <= 'd3; 4914: data <= 'd5; 4915: data <= 'd5; 4916: data <= 'd3; 4917: data <= 'd3; 4918: data <= 'd1; 4919: data <= 'd2; 4920: data <= 'd0; 4921: data <= 'd0; 4922: data <= 'd0; 4923: data <= 'd0; 4924: data <= 'd0; 4925: data <= 'd0; 4926: data <= 'd0; 4927: data <= 'd0; 4928: data <= 'd0; 4929: data <= 'd0; 4930: data <= 'd0; 4931: data <= 'd0; 4932: data <= 'd0; 4933: data <= 'd0; 4934: data <= 'd0; 4935: data <= 'd0; 4936: data <= 'd0; 4937: data <= 'd2; 4938: data <= 'd7; 4939: data <= 'd7; 4940: data <= 'd7; 4941: data <= 'd1; 4942: data <= 'd1; 4943: data <= 'd3; 4944: data <= 'd3; 4945: data <= 'd3; 4946: data <= 'd1; 4947: data <= 'd1; 4948: data <= 'd3; 4949: data <= 'd3; 4950: data <= 'd1; 4951: data <= 'd2; 4952: data <= 'd0; 4953: data <= 'd0; 4954: data <= 'd0; 4955: data <= 'd0; 4956: data <= 'd0; 4957: data <= 'd0; 4958: data <= 'd0; 4959: data <= 'd0; 4960: data <= 'd0; 4961: data <= 'd0; 4962: data <= 'd0; 4963: data <= 'd0; 4964: data <= 'd0; 4965: data <= 'd0; 4966: data <= 'd0; 4967: data <= 'd0; 4968: data <= 'd2; 4969: data <= 'd8; 4970: data <= 'd10; 4971: data <= 'd10; 4972: data <= 'd5; 4973: data <= 'd1; 4974: data <= 'd1; 4975: data <= 'd1; 4976: data <= 'd3; 4977: data <= 'd3; 4978: data <= 'd1; 4979: data <= 'd1; 4980: data <= 'd3; 4981: data <= 'd1; 4982: data <= 'd1; 4983: data <= 'd2; 4984: data <= 'd0; 4985: data <= 'd0; 4986: data <= 'd0; 4987: data <= 'd0; 4988: data <= 'd0; 4989: data <= 'd0; 4990: data <= 'd0; 4991: data <= 'd0; 4992: data <= 'd0; 4993: data <= 'd0; 4994: data <= 'd0; 4995: data <= 'd0; 4996: data <= 'd0; 4997: data <= 'd0; 4998: data <= 'd0; 4999: data <= 'd0; 5000: data <= 'd2; 5001: data <= 'd9; 5002: data <= 'd10; 5003: data <= 'd9; 5004: data <= 'd2; 5005: data <= 'd2; 5006: data <= 'd2; 5007: data <= 'd2; 5008: data <= 'd2; 5009: data <= 'd5; 5010: data <= 'd5; 5011: data <= 'd5; 5012: data <= 'd2; 5013: data <= 'd2; 5014: data <= 'd2; 5015: data <= 'd2; 5016: data <= 'd0; 5017: data <= 'd0; 5018: data <= 'd0; 5019: data <= 'd0; 5020: data <= 'd0; 5021: data <= 'd0; 5022: data <= 'd0; 5023: data <= 'd0; 5024: data <= 'd0; 5025: data <= 'd0; 5026: data <= 'd0; 5027: data <= 'd0; 5028: data <= 'd0; 5029: data <= 'd0; 5030: data <= 'd0; 5031: data <= 'd0; 5032: data <= 'd0; 5033: data <= 'd2; 5034: data <= 'd2; 5035: data <= 'd2; 5036: data <= 'd2; 5037: data <= 'd1; 5038: data <= 'd1; 5039: data <= 'd3; 5040: data <= 'd3; 5041: data <= 'd3; 5042: data <= 'd1; 5043: data <= 'd3; 5044: data <= 'd3; 5045: data <= 'd3; 5046: data <= 'd2; 5047: data <= 'd0; 5048: data <= 'd0; 5049: data <= 'd0; 5050: data <= 'd0; 5051: data <= 'd0; 5052: data <= 'd0; 5053: data <= 'd0; 5054: data <= 'd0; 5055: data <= 'd0; 5056: data <= 'd0; 5057: data <= 'd0; 5058: data <= 'd0; 5059: data <= 'd0; 5060: data <= 'd0; 5061: data <= 'd0; 5062: data <= 'd0; 5063: data <= 'd0; 5064: data <= 'd0; 5065: data <= 'd0; 5066: data <= 'd0; 5067: data <= 'd0; 5068: data <= 'd2; 5069: data <= 'd4; 5070: data <= 'd7; 5071: data <= 'd7; 5072: data <= 'd2; 5073: data <= 'd2; 5074: data <= 'd2; 5075: data <= 'd5; 5076: data <= 'd5; 5077: data <= 'd4; 5078: data <= 'd2; 5079: data <= 'd0; 5080: data <= 'd0; 5081: data <= 'd0; 5082: data <= 'd0; 5083: data <= 'd0; 5084: data <= 'd0; 5085: data <= 'd0; 5086: data <= 'd0; 5087: data <= 'd0; 5088: data <= 'd0; 5089: data <= 'd0; 5090: data <= 'd0; 5091: data <= 'd0; 5092: data <= 'd0; 5093: data <= 'd0; 5094: data <= 'd0; 5095: data <= 'd0; 5096: data <= 'd0; 5097: data <= 'd0; 5098: data <= 'd0; 5099: data <= 'd0; 5100: data <= 'd0; 5101: data <= 'd2; 5102: data <= 'd2; 5103: data <= 'd2; 5104: data <= 'd0; 5105: data <= 'd0; 5106: data <= 'd0; 5107: data <= 'd2; 5108: data <= 'd2; 5109: data <= 'd2; 5110: data <= 'd0; 5111: data <= 'd0; 5112: data <= 'd0; 5113: data <= 'd0; 5114: data <= 'd0; 5115: data <= 'd0; 5116: data <= 'd0; 5117: data <= 'd0; 5118: data <= 'd0; 5119: data <= 'd0; 5120: data <= 'd0; 5121: data <= 'd0; 5122: data <= 'd0; 5123: data <= 'd0; 5124: data <= 'd0; 5125: data <= 'd0; 5126: data <= 'd0; 5127: data <= 'd0; 5128: data <= 'd0; 5129: data <= 'd0; 5130: data <= 'd0; 5131: data <= 'd0; 5132: data <= 'd0; 5133: data <= 'd0; 5134: data <= 'd0; 5135: data <= 'd0; 5136: data <= 'd0; 5137: data <= 'd0; 5138: data <= 'd0; 5139: data <= 'd0; 5140: data <= 'd0; 5141: data <= 'd0; 5142: data <= 'd0; 5143: data <= 'd0; 5144: data <= 'd0; 5145: data <= 'd0; 5146: data <= 'd0; 5147: data <= 'd0; 5148: data <= 'd0; 5149: data <= 'd0; 5150: data <= 'd0; 5151: data <= 'd0; 5152: data <= 'd0; 5153: data <= 'd0; 5154: data <= 'd0; 5155: data <= 'd0; 5156: data <= 'd0; 5157: data <= 'd0; 5158: data <= 'd0; 5159: data <= 'd0; 5160: data <= 'd0; 5161: data <= 'd0; 5162: data <= 'd0; 5163: data <= 'd0; 5164: data <= 'd0; 5165: data <= 'd0; 5166: data <= 'd0; 5167: data <= 'd0; 5168: data <= 'd0; 5169: data <= 'd0; 5170: data <= 'd0; 5171: data <= 'd0; 5172: data <= 'd0; 5173: data <= 'd0; 5174: data <= 'd0; 5175: data <= 'd0; 5176: data <= 'd0; 5177: data <= 'd0; 5178: data <= 'd0; 5179: data <= 'd0; 5180: data <= 'd0; 5181: data <= 'd0; 5182: data <= 'd0; 5183: data <= 'd0; 5184: data <= 'd0; 5185: data <= 'd0; 5186: data <= 'd0; 5187: data <= 'd0; 5188: data <= 'd0; 5189: data <= 'd0; 5190: data <= 'd0; 5191: data <= 'd0; 5192: data <= 'd0; 5193: data <= 'd0; 5194: data <= 'd0; 5195: data <= 'd0; 5196: data <= 'd0; 5197: data <= 'd0; 5198: data <= 'd0; 5199: data <= 'd0; 5200: data <= 'd0; 5201: data <= 'd0; 5202: data <= 'd0; 5203: data <= 'd0; 5204: data <= 'd0; 5205: data <= 'd0; 5206: data <= 'd0; 5207: data <= 'd0; 5208: data <= 'd0; 5209: data <= 'd0; 5210: data <= 'd0; 5211: data <= 'd0; 5212: data <= 'd0; 5213: data <= 'd0; 5214: data <= 'd0; 5215: data <= 'd0; 5216: data <= 'd0; 5217: data <= 'd0; 5218: data <= 'd0; 5219: data <= 'd0; 5220: data <= 'd0; 5221: data <= 'd0; 5222: data <= 'd0; 5223: data <= 'd0; 5224: data <= 'd0; 5225: data <= 'd0; 5226: data <= 'd0; 5227: data <= 'd0; 5228: data <= 'd0; 5229: data <= 'd0; 5230: data <= 'd0; 5231: data <= 'd0; 5232: data <= 'd0; 5233: data <= 'd0; 5234: data <= 'd0; 5235: data <= 'd0; 5236: data <= 'd0; 5237: data <= 'd0; 5238: data <= 'd0; 5239: data <= 'd0; 5240: data <= 'd0; 5241: data <= 'd0; 5242: data <= 'd0; 5243: data <= 'd0; 5244: data <= 'd0; 5245: data <= 'd0; 5246: data <= 'd0; 5247: data <= 'd0; 5248: data <= 'd0; 5249: data <= 'd0; 5250: data <= 'd0; 5251: data <= 'd0; 5252: data <= 'd0; 5253: data <= 'd0; 5254: data <= 'd0; 5255: data <= 'd0; 5256: data <= 'd0; 5257: data <= 'd0; 5258: data <= 'd0; 5259: data <= 'd0; 5260: data <= 'd0; 5261: data <= 'd0; 5262: data <= 'd0; 5263: data <= 'd0; 5264: data <= 'd0; 5265: data <= 'd0; 5266: data <= 'd0; 5267: data <= 'd0; 5268: data <= 'd0; 5269: data <= 'd0; 5270: data <= 'd0; 5271: data <= 'd0; 5272: data <= 'd0; 5273: data <= 'd0; 5274: data <= 'd0; 5275: data <= 'd0; 5276: data <= 'd0; 5277: data <= 'd0; 5278: data <= 'd0; 5279: data <= 'd0; 5280: data <= 'd0; 5281: data <= 'd0; 5282: data <= 'd0; 5283: data <= 'd0; 5284: data <= 'd0; 5285: data <= 'd0; 5286: data <= 'd0; 5287: data <= 'd0; 5288: data <= 'd0; 5289: data <= 'd0; 5290: data <= 'd0; 5291: data <= 'd0; 5292: data <= 'd0; 5293: data <= 'd0; 5294: data <= 'd0; 5295: data <= 'd0; 5296: data <= 'd0; 5297: data <= 'd0; 5298: data <= 'd0; 5299: data <= 'd0; 5300: data <= 'd0; 5301: data <= 'd0; 5302: data <= 'd0; 5303: data <= 'd0; 5304: data <= 'd0; 5305: data <= 'd0; 5306: data <= 'd0; 5307: data <= 'd0; 5308: data <= 'd0; 5309: data <= 'd0; 5310: data <= 'd0; 5311: data <= 'd0; 5312: data <= 'd0; 5313: data <= 'd0; 5314: data <= 'd0; 5315: data <= 'd0; 5316: data <= 'd0; 5317: data <= 'd0; 5318: data <= 'd0; 5319: data <= 'd0; 5320: data <= 'd0; 5321: data <= 'd0; 5322: data <= 'd0; 5323: data <= 'd0; 5324: data <= 'd0; 5325: data <= 'd0; 5326: data <= 'd0; 5327: data <= 'd0; 5328: data <= 'd0; 5329: data <= 'd0; 5330: data <= 'd0; 5331: data <= 'd0; 5332: data <= 'd0; 5333: data <= 'd0; 5334: data <= 'd0; 5335: data <= 'd0; 5336: data <= 'd0; 5337: data <= 'd0; 5338: data <= 'd0; 5339: data <= 'd0; 5340: data <= 'd0; 5341: data <= 'd0; 5342: data <= 'd0; 5343: data <= 'd0; 5344: data <= 'd0; 5345: data <= 'd0; 5346: data <= 'd0; 5347: data <= 'd0; 5348: data <= 'd0; 5349: data <= 'd0; 5350: data <= 'd0; 5351: data <= 'd0; 5352: data <= 'd0; 5353: data <= 'd0; 5354: data <= 'd0; 5355: data <= 'd0; 5356: data <= 'd0; 5357: data <= 'd0; 5358: data <= 'd0; 5359: data <= 'd0; 5360: data <= 'd0; 5361: data <= 'd0; 5362: data <= 'd0; 5363: data <= 'd0; 5364: data <= 'd0; 5365: data <= 'd0; 5366: data <= 'd0; 5367: data <= 'd0; 5368: data <= 'd0; 5369: data <= 'd0; 5370: data <= 'd0; 5371: data <= 'd0; 5372: data <= 'd0; 5373: data <= 'd0; 5374: data <= 'd0; 5375: data <= 'd0; 5376: data <= 'd0; 5377: data <= 'd0; 5378: data <= 'd0; 5379: data <= 'd0; 5380: data <= 'd0; 5381: data <= 'd0; 5382: data <= 'd0; 5383: data <= 'd0; 5384: data <= 'd0; 5385: data <= 'd0; 5386: data <= 'd0; 5387: data <= 'd0; 5388: data <= 'd0; 5389: data <= 'd2; 5390: data <= 'd2; 5391: data <= 'd2; 5392: data <= 'd2; 5393: data <= 'd2; 5394: data <= 'd2; 5395: data <= 'd0; 5396: data <= 'd0; 5397: data <= 'd0; 5398: data <= 'd0; 5399: data <= 'd0; 5400: data <= 'd0; 5401: data <= 'd0; 5402: data <= 'd0; 5403: data <= 'd0; 5404: data <= 'd0; 5405: data <= 'd0; 5406: data <= 'd0; 5407: data <= 'd0; 5408: data <= 'd0; 5409: data <= 'd0; 5410: data <= 'd0; 5411: data <= 'd0; 5412: data <= 'd0; 5413: data <= 'd0; 5414: data <= 'd0; 5415: data <= 'd0; 5416: data <= 'd0; 5417: data <= 'd0; 5418: data <= 'd0; 5419: data <= 'd2; 5420: data <= 'd2; 5421: data <= 'd6; 5422: data <= 'd6; 5423: data <= 'd6; 5424: data <= 'd6; 5425: data <= 'd6; 5426: data <= 'd6; 5427: data <= 'd2; 5428: data <= 'd2; 5429: data <= 'd0; 5430: data <= 'd0; 5431: data <= 'd0; 5432: data <= 'd0; 5433: data <= 'd0; 5434: data <= 'd0; 5435: data <= 'd0; 5436: data <= 'd0; 5437: data <= 'd0; 5438: data <= 'd0; 5439: data <= 'd0; 5440: data <= 'd0; 5441: data <= 'd0; 5442: data <= 'd0; 5443: data <= 'd0; 5444: data <= 'd0; 5445: data <= 'd0; 5446: data <= 'd0; 5447: data <= 'd0; 5448: data <= 'd0; 5449: data <= 'd0; 5450: data <= 'd2; 5451: data <= 'd1; 5452: data <= 'd3; 5453: data <= 'd6; 5454: data <= 'd6; 5455: data <= 'd6; 5456: data <= 'd6; 5457: data <= 'd6; 5458: data <= 'd6; 5459: data <= 'd6; 5460: data <= 'd3; 5461: data <= 'd2; 5462: data <= 'd0; 5463: data <= 'd0; 5464: data <= 'd0; 5465: data <= 'd0; 5466: data <= 'd0; 5467: data <= 'd0; 5468: data <= 'd0; 5469: data <= 'd0; 5470: data <= 'd0; 5471: data <= 'd0; 5472: data <= 'd0; 5473: data <= 'd0; 5474: data <= 'd0; 5475: data <= 'd0; 5476: data <= 'd0; 5477: data <= 'd0; 5478: data <= 'd0; 5479: data <= 'd0; 5480: data <= 'd0; 5481: data <= 'd2; 5482: data <= 'd1; 5483: data <= 'd1; 5484: data <= 'd1; 5485: data <= 'd3; 5486: data <= 'd6; 5487: data <= 'd6; 5488: data <= 'd6; 5489: data <= 'd6; 5490: data <= 'd6; 5491: data <= 'd3; 5492: data <= 'd1; 5493: data <= 'd1; 5494: data <= 'd2; 5495: data <= 'd0; 5496: data <= 'd0; 5497: data <= 'd0; 5498: data <= 'd0; 5499: data <= 'd0; 5500: data <= 'd0; 5501: data <= 'd0; 5502: data <= 'd0; 5503: data <= 'd0; 5504: data <= 'd0; 5505: data <= 'd0; 5506: data <= 'd0; 5507: data <= 'd0; 5508: data <= 'd0; 5509: data <= 'd0; 5510: data <= 'd0; 5511: data <= 'd0; 5512: data <= 'd0; 5513: data <= 'd2; 5514: data <= 'd1; 5515: data <= 'd1; 5516: data <= 'd5; 5517: data <= 'd5; 5518: data <= 'd5; 5519: data <= 'd1; 5520: data <= 'd1; 5521: data <= 'd1; 5522: data <= 'd1; 5523: data <= 'd1; 5524: data <= 'd5; 5525: data <= 'd5; 5526: data <= 'd2; 5527: data <= 'd0; 5528: data <= 'd0; 5529: data <= 'd0; 5530: data <= 'd0; 5531: data <= 'd0; 5532: data <= 'd0; 5533: data <= 'd0; 5534: data <= 'd0; 5535: data <= 'd0; 5536: data <= 'd0; 5537: data <= 'd0; 5538: data <= 'd0; 5539: data <= 'd0; 5540: data <= 'd0; 5541: data <= 'd0; 5542: data <= 'd0; 5543: data <= 'd0; 5544: data <= 'd2; 5545: data <= 'd1; 5546: data <= 'd5; 5547: data <= 'd5; 5548: data <= 'd3; 5549: data <= 'd6; 5550: data <= 'd6; 5551: data <= 'd6; 5552: data <= 'd6; 5553: data <= 'd6; 5554: data <= 'd6; 5555: data <= 'd6; 5556: data <= 'd6; 5557: data <= 'd3; 5558: data <= 'd5; 5559: data <= 'd2; 5560: data <= 'd0; 5561: data <= 'd0; 5562: data <= 'd0; 5563: data <= 'd0; 5564: data <= 'd0; 5565: data <= 'd0; 5566: data <= 'd0; 5567: data <= 'd0; 5568: data <= 'd0; 5569: data <= 'd0; 5570: data <= 'd0; 5571: data <= 'd0; 5572: data <= 'd0; 5573: data <= 'd0; 5574: data <= 'd0; 5575: data <= 'd0; 5576: data <= 'd2; 5577: data <= 'd5; 5578: data <= 'd3; 5579: data <= 'd6; 5580: data <= 'd3; 5581: data <= 'd1; 5582: data <= 'd1; 5583: data <= 'd1; 5584: data <= 'd1; 5585: data <= 'd1; 5586: data <= 'd1; 5587: data <= 'd1; 5588: data <= 'd1; 5589: data <= 'd1; 5590: data <= 'd3; 5591: data <= 'd2; 5592: data <= 'd0; 5593: data <= 'd0; 5594: data <= 'd0; 5595: data <= 'd0; 5596: data <= 'd0; 5597: data <= 'd0; 5598: data <= 'd0; 5599: data <= 'd0; 5600: data <= 'd0; 5601: data <= 'd0; 5602: data <= 'd0; 5603: data <= 'd0; 5604: data <= 'd0; 5605: data <= 'd0; 5606: data <= 'd0; 5607: data <= 'd0; 5608: data <= 'd2; 5609: data <= 'd5; 5610: data <= 'd3; 5611: data <= 'd1; 5612: data <= 'd1; 5613: data <= 'd1; 5614: data <= 'd5; 5615: data <= 'd5; 5616: data <= 'd5; 5617: data <= 'd5; 5618: data <= 'd5; 5619: data <= 'd5; 5620: data <= 'd5; 5621: data <= 'd1; 5622: data <= 'd1; 5623: data <= 'd2; 5624: data <= 'd0; 5625: data <= 'd0; 5626: data <= 'd0; 5627: data <= 'd0; 5628: data <= 'd0; 5629: data <= 'd0; 5630: data <= 'd0; 5631: data <= 'd0; 5632: data <= 'd0; 5633: data <= 'd0; 5634: data <= 'd0; 5635: data <= 'd0; 5636: data <= 'd0; 5637: data <= 'd0; 5638: data <= 'd0; 5639: data <= 'd0; 5640: data <= 'd2; 5641: data <= 'd6; 5642: data <= 'd1; 5643: data <= 'd5; 5644: data <= 'd2; 5645: data <= 'd2; 5646: data <= 'd2; 5647: data <= 'd2; 5648: data <= 'd2; 5649: data <= 'd2; 5650: data <= 'd2; 5651: data <= 'd2; 5652: data <= 'd2; 5653: data <= 'd2; 5654: data <= 'd5; 5655: data <= 'd2; 5656: data <= 'd0; 5657: data <= 'd0; 5658: data <= 'd0; 5659: data <= 'd0; 5660: data <= 'd0; 5661: data <= 'd0; 5662: data <= 'd0; 5663: data <= 'd0; 5664: data <= 'd0; 5665: data <= 'd0; 5666: data <= 'd0; 5667: data <= 'd0; 5668: data <= 'd0; 5669: data <= 'd0; 5670: data <= 'd0; 5671: data <= 'd0; 5672: data <= 'd2; 5673: data <= 'd1; 5674: data <= 'd5; 5675: data <= 'd2; 5676: data <= 'd8; 5677: data <= 'd8; 5678: data <= 'd8; 5679: data <= 'd8; 5680: data <= 'd8; 5681: data <= 'd9; 5682: data <= 'd9; 5683: data <= 'd8; 5684: data <= 'd8; 5685: data <= 'd8; 5686: data <= 'd2; 5687: data <= 'd2; 5688: data <= 'd0; 5689: data <= 'd0; 5690: data <= 'd0; 5691: data <= 'd0; 5692: data <= 'd0; 5693: data <= 'd0; 5694: data <= 'd0; 5695: data <= 'd0; 5696: data <= 'd0; 5697: data <= 'd0; 5698: data <= 'd0; 5699: data <= 'd0; 5700: data <= 'd0; 5701: data <= 'd0; 5702: data <= 'd2; 5703: data <= 'd2; 5704: data <= 'd2; 5705: data <= 'd1; 5706: data <= 'd2; 5707: data <= 'd8; 5708: data <= 'd8; 5709: data <= 'd9; 5710: data <= 'd9; 5711: data <= 'd2; 5712: data <= 'd9; 5713: data <= 'd11; 5714: data <= 'd11; 5715: data <= 'd10; 5716: data <= 'd2; 5717: data <= 'd9; 5718: data <= 'd2; 5719: data <= 'd2; 5720: data <= 'd0; 5721: data <= 'd0; 5722: data <= 'd0; 5723: data <= 'd0; 5724: data <= 'd0; 5725: data <= 'd0; 5726: data <= 'd0; 5727: data <= 'd0; 5728: data <= 'd0; 5729: data <= 'd0; 5730: data <= 'd0; 5731: data <= 'd0; 5732: data <= 'd0; 5733: data <= 'd0; 5734: data <= 'd2; 5735: data <= 'd1; 5736: data <= 'd1; 5737: data <= 'd2; 5738: data <= 'd9; 5739: data <= 'd10; 5740: data <= 'd9; 5741: data <= 'd9; 5742: data <= 'd10; 5743: data <= 'd11; 5744: data <= 'd10; 5745: data <= 'd11; 5746: data <= 'd11; 5747: data <= 'd10; 5748: data <= 'd11; 5749: data <= 'd10; 5750: data <= 'd9; 5751: data <= 'd2; 5752: data <= 'd0; 5753: data <= 'd0; 5754: data <= 'd0; 5755: data <= 'd0; 5756: data <= 'd0; 5757: data <= 'd0; 5758: data <= 'd0; 5759: data <= 'd0; 5760: data <= 'd0; 5761: data <= 'd0; 5762: data <= 'd0; 5763: data <= 'd0; 5764: data <= 'd0; 5765: data <= 'd0; 5766: data <= 'd2; 5767: data <= 'd5; 5768: data <= 'd5; 5769: data <= 'd5; 5770: data <= 'd2; 5771: data <= 'd8; 5772: data <= 'd9; 5773: data <= 'd9; 5774: data <= 'd10; 5775: data <= 'd10; 5776: data <= 'd10; 5777: data <= 'd8; 5778: data <= 'd8; 5779: data <= 'd10; 5780: data <= 'd10; 5781: data <= 'd9; 5782: data <= 'd2; 5783: data <= 'd0; 5784: data <= 'd0; 5785: data <= 'd0; 5786: data <= 'd0; 5787: data <= 'd0; 5788: data <= 'd0; 5789: data <= 'd0; 5790: data <= 'd0; 5791: data <= 'd0; 5792: data <= 'd0; 5793: data <= 'd0; 5794: data <= 'd0; 5795: data <= 'd0; 5796: data <= 'd0; 5797: data <= 'd0; 5798: data <= 'd0; 5799: data <= 'd2; 5800: data <= 'd2; 5801: data <= 'd2; 5802: data <= 'd2; 5803: data <= 'd8; 5804: data <= 'd8; 5805: data <= 'd9; 5806: data <= 'd9; 5807: data <= 'd10; 5808: data <= 'd10; 5809: data <= 'd9; 5810: data <= 'd9; 5811: data <= 'd10; 5812: data <= 'd10; 5813: data <= 'd9; 5814: data <= 'd2; 5815: data <= 'd0; 5816: data <= 'd0; 5817: data <= 'd0; 5818: data <= 'd0; 5819: data <= 'd0; 5820: data <= 'd0; 5821: data <= 'd0; 5822: data <= 'd0; 5823: data <= 'd0; 5824: data <= 'd0; 5825: data <= 'd0; 5826: data <= 'd0; 5827: data <= 'd0; 5828: data <= 'd0; 5829: data <= 'd0; 5830: data <= 'd0; 5831: data <= 'd0; 5832: data <= 'd0; 5833: data <= 'd0; 5834: data <= 'd2; 5835: data <= 'd2; 5836: data <= 'd5; 5837: data <= 'd5; 5838: data <= 'd8; 5839: data <= 'd9; 5840: data <= 'd9; 5841: data <= 'd9; 5842: data <= 'd9; 5843: data <= 'd9; 5844: data <= 'd9; 5845: data <= 'd5; 5846: data <= 'd2; 5847: data <= 'd0; 5848: data <= 'd0; 5849: data <= 'd0; 5850: data <= 'd0; 5851: data <= 'd0; 5852: data <= 'd0; 5853: data <= 'd0; 5854: data <= 'd0; 5855: data <= 'd0; 5856: data <= 'd0; 5857: data <= 'd0; 5858: data <= 'd0; 5859: data <= 'd0; 5860: data <= 'd0; 5861: data <= 'd0; 5862: data <= 'd0; 5863: data <= 'd0; 5864: data <= 'd0; 5865: data <= 'd2; 5866: data <= 'd7; 5867: data <= 'd1; 5868: data <= 'd1; 5869: data <= 'd1; 5870: data <= 'd3; 5871: data <= 'd3; 5872: data <= 'd3; 5873: data <= 'd5; 5874: data <= 'd5; 5875: data <= 'd3; 5876: data <= 'd3; 5877: data <= 'd1; 5878: data <= 'd2; 5879: data <= 'd0; 5880: data <= 'd0; 5881: data <= 'd0; 5882: data <= 'd0; 5883: data <= 'd0; 5884: data <= 'd0; 5885: data <= 'd0; 5886: data <= 'd0; 5887: data <= 'd0; 5888: data <= 'd0; 5889: data <= 'd0; 5890: data <= 'd0; 5891: data <= 'd0; 5892: data <= 'd0; 5893: data <= 'd0; 5894: data <= 'd0; 5895: data <= 'd0; 5896: data <= 'd0; 5897: data <= 'd2; 5898: data <= 'd7; 5899: data <= 'd7; 5900: data <= 'd1; 5901: data <= 'd1; 5902: data <= 'd3; 5903: data <= 'd3; 5904: data <= 'd3; 5905: data <= 'd1; 5906: data <= 'd1; 5907: data <= 'd3; 5908: data <= 'd3; 5909: data <= 'd1; 5910: data <= 'd2; 5911: data <= 'd0; 5912: data <= 'd0; 5913: data <= 'd0; 5914: data <= 'd0; 5915: data <= 'd0; 5916: data <= 'd0; 5917: data <= 'd0; 5918: data <= 'd0; 5919: data <= 'd0; 5920: data <= 'd0; 5921: data <= 'd0; 5922: data <= 'd0; 5923: data <= 'd0; 5924: data <= 'd0; 5925: data <= 'd0; 5926: data <= 'd0; 5927: data <= 'd0; 5928: data <= 'd2; 5929: data <= 'd9; 5930: data <= 'd9; 5931: data <= 'd7; 5932: data <= 'd1; 5933: data <= 'd1; 5934: data <= 'd1; 5935: data <= 'd3; 5936: data <= 'd3; 5937: data <= 'd1; 5938: data <= 'd1; 5939: data <= 'd3; 5940: data <= 'd1; 5941: data <= 'd1; 5942: data <= 'd8; 5943: data <= 'd2; 5944: data <= 'd0; 5945: data <= 'd0; 5946: data <= 'd0; 5947: data <= 'd0; 5948: data <= 'd0; 5949: data <= 'd0; 5950: data <= 'd0; 5951: data <= 'd0; 5952: data <= 'd0; 5953: data <= 'd0; 5954: data <= 'd0; 5955: data <= 'd0; 5956: data <= 'd0; 5957: data <= 'd0; 5958: data <= 'd0; 5959: data <= 'd0; 5960: data <= 'd2; 5961: data <= 'd9; 5962: data <= 'd9; 5963: data <= 'd2; 5964: data <= 'd2; 5965: data <= 'd2; 5966: data <= 'd2; 5967: data <= 'd2; 5968: data <= 'd5; 5969: data <= 'd5; 5970: data <= 'd5; 5971: data <= 'd2; 5972: data <= 'd2; 5973: data <= 'd2; 5974: data <= 'd8; 5975: data <= 'd2; 5976: data <= 'd0; 5977: data <= 'd0; 5978: data <= 'd0; 5979: data <= 'd0; 5980: data <= 'd0; 5981: data <= 'd0; 5982: data <= 'd0; 5983: data <= 'd0; 5984: data <= 'd0; 5985: data <= 'd0; 5986: data <= 'd0; 5987: data <= 'd0; 5988: data <= 'd0; 5989: data <= 'd0; 5990: data <= 'd0; 5991: data <= 'd0; 5992: data <= 'd0; 5993: data <= 'd2; 5994: data <= 'd2; 5995: data <= 'd2; 5996: data <= 'd1; 5997: data <= 'd1; 5998: data <= 'd3; 5999: data <= 'd3; 6000: data <= 'd3; 6001: data <= 'd1; 6002: data <= 'd3; 6003: data <= 'd3; 6004: data <= 'd3; 6005: data <= 'd2; 6006: data <= 'd2; 6007: data <= 'd0; 6008: data <= 'd0; 6009: data <= 'd0; 6010: data <= 'd0; 6011: data <= 'd0; 6012: data <= 'd0; 6013: data <= 'd0; 6014: data <= 'd0; 6015: data <= 'd0; 6016: data <= 'd0; 6017: data <= 'd0; 6018: data <= 'd0; 6019: data <= 'd0; 6020: data <= 'd0; 6021: data <= 'd0; 6022: data <= 'd0; 6023: data <= 'd0; 6024: data <= 'd0; 6025: data <= 'd0; 6026: data <= 'd0; 6027: data <= 'd2; 6028: data <= 'd4; 6029: data <= 'd7; 6030: data <= 'd7; 6031: data <= 'd2; 6032: data <= 'd2; 6033: data <= 'd2; 6034: data <= 'd5; 6035: data <= 'd5; 6036: data <= 'd4; 6037: data <= 'd2; 6038: data <= 'd0; 6039: data <= 'd0; 6040: data <= 'd0; 6041: data <= 'd0; 6042: data <= 'd0; 6043: data <= 'd0; 6044: data <= 'd0; 6045: data <= 'd0; 6046: data <= 'd0; 6047: data <= 'd0; 6048: data <= 'd0; 6049: data <= 'd0; 6050: data <= 'd0; 6051: data <= 'd0; 6052: data <= 'd0; 6053: data <= 'd0; 6054: data <= 'd0; 6055: data <= 'd0; 6056: data <= 'd0; 6057: data <= 'd0; 6058: data <= 'd0; 6059: data <= 'd2; 6060: data <= 'd4; 6061: data <= 'd7; 6062: data <= 'd2; 6063: data <= 'd0; 6064: data <= 'd0; 6065: data <= 'd0; 6066: data <= 'd2; 6067: data <= 'd4; 6068: data <= 'd4; 6069: data <= 'd2; 6070: data <= 'd0; 6071: data <= 'd0; 6072: data <= 'd0; 6073: data <= 'd0; 6074: data <= 'd0; 6075: data <= 'd0; 6076: data <= 'd0; 6077: data <= 'd0; 6078: data <= 'd0; 6079: data <= 'd0; 6080: data <= 'd0; 6081: data <= 'd0; 6082: data <= 'd0; 6083: data <= 'd0; 6084: data <= 'd0; 6085: data <= 'd0; 6086: data <= 'd0; 6087: data <= 'd0; 6088: data <= 'd0; 6089: data <= 'd0; 6090: data <= 'd0; 6091: data <= 'd2; 6092: data <= 'd2; 6093: data <= 'd2; 6094: data <= 'd0; 6095: data <= 'd0; 6096: data <= 'd0; 6097: data <= 'd0; 6098: data <= 'd2; 6099: data <= 'd2; 6100: data <= 'd2; 6101: data <= 'd0; 6102: data <= 'd0; 6103: data <= 'd0; 6104: data <= 'd0; 6105: data <= 'd0; 6106: data <= 'd0; 6107: data <= 'd0; 6108: data <= 'd0; 6109: data <= 'd0; 6110: data <= 'd0; 6111: data <= 'd0; 6112: data <= 'd0; 6113: data <= 'd0; 6114: data <= 'd0; 6115: data <= 'd0; 6116: data <= 'd0; 6117: data <= 'd0; 6118: data <= 'd0; 6119: data <= 'd0; 6120: data <= 'd0; 6121: data <= 'd0; 6122: data <= 'd0; 6123: data <= 'd0; 6124: data <= 'd0; 6125: data <= 'd0; 6126: data <= 'd0; 6127: data <= 'd0; 6128: data <= 'd0; 6129: data <= 'd0; 6130: data <= 'd0; 6131: data <= 'd0; 6132: data <= 'd0; 6133: data <= 'd0; 6134: data <= 'd0; 6135: data <= 'd0; 6136: data <= 'd0; 6137: data <= 'd0; 6138: data <= 'd0; 6139: data <= 'd0; 6140: data <= 'd0; 6141: data <= 'd0; 6142: data <= 'd0; 6143: data <= 'd0; 6144: data <= 'd0; 6145: data <= 'd0; 6146: data <= 'd0; 6147: data <= 'd0; 6148: data <= 'd0; 6149: data <= 'd0; 6150: data <= 'd0; 6151: data <= 'd0; 6152: data <= 'd0; 6153: data <= 'd0; 6154: data <= 'd0; 6155: data <= 'd0; 6156: data <= 'd0; 6157: data <= 'd0; 6158: data <= 'd0; 6159: data <= 'd0; 6160: data <= 'd0; 6161: data <= 'd0; 6162: data <= 'd0; 6163: data <= 'd0; 6164: data <= 'd0; 6165: data <= 'd0; 6166: data <= 'd0; 6167: data <= 'd0; 6168: data <= 'd0; 6169: data <= 'd0; 6170: data <= 'd0; 6171: data <= 'd0; 6172: data <= 'd0; 6173: data <= 'd0; 6174: data <= 'd0; 6175: data <= 'd0; 6176: data <= 'd0; 6177: data <= 'd0; 6178: data <= 'd0; 6179: data <= 'd0; 6180: data <= 'd0; 6181: data <= 'd0; 6182: data <= 'd0; 6183: data <= 'd0; 6184: data <= 'd0; 6185: data <= 'd0; 6186: data <= 'd0; 6187: data <= 'd0; 6188: data <= 'd0; 6189: data <= 'd0; 6190: data <= 'd0; 6191: data <= 'd0; 6192: data <= 'd0; 6193: data <= 'd0; 6194: data <= 'd0; 6195: data <= 'd0; 6196: data <= 'd0; 6197: data <= 'd0; 6198: data <= 'd0; 6199: data <= 'd0; 6200: data <= 'd0; 6201: data <= 'd0; 6202: data <= 'd0; 6203: data <= 'd0; 6204: data <= 'd0; 6205: data <= 'd0; 6206: data <= 'd0; 6207: data <= 'd0; 6208: data <= 'd0; 6209: data <= 'd0; 6210: data <= 'd0; 6211: data <= 'd0; 6212: data <= 'd0; 6213: data <= 'd0; 6214: data <= 'd0; 6215: data <= 'd0; 6216: data <= 'd0; 6217: data <= 'd0; 6218: data <= 'd0; 6219: data <= 'd0; 6220: data <= 'd0; 6221: data <= 'd0; 6222: data <= 'd0; 6223: data <= 'd0; 6224: data <= 'd0; 6225: data <= 'd0; 6226: data <= 'd0; 6227: data <= 'd0; 6228: data <= 'd0; 6229: data <= 'd0; 6230: data <= 'd0; 6231: data <= 'd0; 6232: data <= 'd0; 6233: data <= 'd0; 6234: data <= 'd0; 6235: data <= 'd0; 6236: data <= 'd0; 6237: data <= 'd0; 6238: data <= 'd0; 6239: data <= 'd0; 6240: data <= 'd0; 6241: data <= 'd0; 6242: data <= 'd0; 6243: data <= 'd0; 6244: data <= 'd0; 6245: data <= 'd0; 6246: data <= 'd0; 6247: data <= 'd0; 6248: data <= 'd0; 6249: data <= 'd0; 6250: data <= 'd0; 6251: data <= 'd0; 6252: data <= 'd0; 6253: data <= 'd0; 6254: data <= 'd0; 6255: data <= 'd0; 6256: data <= 'd0; 6257: data <= 'd0; 6258: data <= 'd0; 6259: data <= 'd0; 6260: data <= 'd0; 6261: data <= 'd0; 6262: data <= 'd0; 6263: data <= 'd0; 6264: data <= 'd0; 6265: data <= 'd0; 6266: data <= 'd0; 6267: data <= 'd0; 6268: data <= 'd0; 6269: data <= 'd0; 6270: data <= 'd0; 6271: data <= 'd0; 6272: data <= 'd0; 6273: data <= 'd0; 6274: data <= 'd0; 6275: data <= 'd0; 6276: data <= 'd0; 6277: data <= 'd0; 6278: data <= 'd0; 6279: data <= 'd0; 6280: data <= 'd0; 6281: data <= 'd0; 6282: data <= 'd0; 6283: data <= 'd0; 6284: data <= 'd0; 6285: data <= 'd0; 6286: data <= 'd0; 6287: data <= 'd0; 6288: data <= 'd0; 6289: data <= 'd0; 6290: data <= 'd0; 6291: data <= 'd0; 6292: data <= 'd0; 6293: data <= 'd0; 6294: data <= 'd0; 6295: data <= 'd0; 6296: data <= 'd0; 6297: data <= 'd0; 6298: data <= 'd0; 6299: data <= 'd0; 6300: data <= 'd0; 6301: data <= 'd0; 6302: data <= 'd0; 6303: data <= 'd0; 6304: data <= 'd0; 6305: data <= 'd0; 6306: data <= 'd0; 6307: data <= 'd0; 6308: data <= 'd0; 6309: data <= 'd0; 6310: data <= 'd0; 6311: data <= 'd0; 6312: data <= 'd0; 6313: data <= 'd0; 6314: data <= 'd0; 6315: data <= 'd0; 6316: data <= 'd0; 6317: data <= 'd0; 6318: data <= 'd0; 6319: data <= 'd0; 6320: data <= 'd0; 6321: data <= 'd0; 6322: data <= 'd0; 6323: data <= 'd0; 6324: data <= 'd0; 6325: data <= 'd0; 6326: data <= 'd0; 6327: data <= 'd0; 6328: data <= 'd0; 6329: data <= 'd0; 6330: data <= 'd0; 6331: data <= 'd0; 6332: data <= 'd0; 6333: data <= 'd0; 6334: data <= 'd0; 6335: data <= 'd0; 6336: data <= 'd0; 6337: data <= 'd0; 6338: data <= 'd0; 6339: data <= 'd0; 6340: data <= 'd0; 6341: data <= 'd0; 6342: data <= 'd0; 6343: data <= 'd0; 6344: data <= 'd0; 6345: data <= 'd0; 6346: data <= 'd0; 6347: data <= 'd0; 6348: data <= 'd0; 6349: data <= 'd0; 6350: data <= 'd0; 6351: data <= 'd0; 6352: data <= 'd0; 6353: data <= 'd0; 6354: data <= 'd0; 6355: data <= 'd0; 6356: data <= 'd0; 6357: data <= 'd0; 6358: data <= 'd0; 6359: data <= 'd0; 6360: data <= 'd0; 6361: data <= 'd0; 6362: data <= 'd0; 6363: data <= 'd0; 6364: data <= 'd0; 6365: data <= 'd0; 6366: data <= 'd0; 6367: data <= 'd0; 6368: data <= 'd0; 6369: data <= 'd0; 6370: data <= 'd0; 6371: data <= 'd0; 6372: data <= 'd0; 6373: data <= 'd0; 6374: data <= 'd0; 6375: data <= 'd0; 6376: data <= 'd0; 6377: data <= 'd0; 6378: data <= 'd0; 6379: data <= 'd0; 6380: data <= 'd0; 6381: data <= 'd0; 6382: data <= 'd0; 6383: data <= 'd0; 6384: data <= 'd0; 6385: data <= 'd0; 6386: data <= 'd0; 6387: data <= 'd0; 6388: data <= 'd0; 6389: data <= 'd0; 6390: data <= 'd0; 6391: data <= 'd0; 6392: data <= 'd0; 6393: data <= 'd0; 6394: data <= 'd0; 6395: data <= 'd0; 6396: data <= 'd0; 6397: data <= 'd0; 6398: data <= 'd0; 6399: data <= 'd0; 6400: data <= 'd0; 6401: data <= 'd0; 6402: data <= 'd0; 6403: data <= 'd0; 6404: data <= 'd0; 6405: data <= 'd0; 6406: data <= 'd0; 6407: data <= 'd0; 6408: data <= 'd0; 6409: data <= 'd0; 6410: data <= 'd0; 6411: data <= 'd0; 6412: data <= 'd0; 6413: data <= 'd2; 6414: data <= 'd2; 6415: data <= 'd2; 6416: data <= 'd2; 6417: data <= 'd2; 6418: data <= 'd2; 6419: data <= 'd0; 6420: data <= 'd0; 6421: data <= 'd0; 6422: data <= 'd0; 6423: data <= 'd0; 6424: data <= 'd0; 6425: data <= 'd0; 6426: data <= 'd0; 6427: data <= 'd0; 6428: data <= 'd0; 6429: data <= 'd0; 6430: data <= 'd0; 6431: data <= 'd0; 6432: data <= 'd0; 6433: data <= 'd0; 6434: data <= 'd0; 6435: data <= 'd0; 6436: data <= 'd0; 6437: data <= 'd0; 6438: data <= 'd0; 6439: data <= 'd0; 6440: data <= 'd0; 6441: data <= 'd0; 6442: data <= 'd0; 6443: data <= 'd2; 6444: data <= 'd2; 6445: data <= 'd6; 6446: data <= 'd6; 6447: data <= 'd6; 6448: data <= 'd6; 6449: data <= 'd6; 6450: data <= 'd6; 6451: data <= 'd2; 6452: data <= 'd2; 6453: data <= 'd0; 6454: data <= 'd0; 6455: data <= 'd0; 6456: data <= 'd0; 6457: data <= 'd0; 6458: data <= 'd0; 6459: data <= 'd0; 6460: data <= 'd0; 6461: data <= 'd0; 6462: data <= 'd0; 6463: data <= 'd0; 6464: data <= 'd0; 6465: data <= 'd0; 6466: data <= 'd0; 6467: data <= 'd0; 6468: data <= 'd0; 6469: data <= 'd0; 6470: data <= 'd0; 6471: data <= 'd0; 6472: data <= 'd0; 6473: data <= 'd0; 6474: data <= 'd2; 6475: data <= 'd1; 6476: data <= 'd3; 6477: data <= 'd6; 6478: data <= 'd6; 6479: data <= 'd6; 6480: data <= 'd6; 6481: data <= 'd6; 6482: data <= 'd6; 6483: data <= 'd6; 6484: data <= 'd3; 6485: data <= 'd2; 6486: data <= 'd0; 6487: data <= 'd0; 6488: data <= 'd0; 6489: data <= 'd0; 6490: data <= 'd0; 6491: data <= 'd0; 6492: data <= 'd0; 6493: data <= 'd0; 6494: data <= 'd0; 6495: data <= 'd0; 6496: data <= 'd0; 6497: data <= 'd0; 6498: data <= 'd0; 6499: data <= 'd0; 6500: data <= 'd0; 6501: data <= 'd0; 6502: data <= 'd0; 6503: data <= 'd0; 6504: data <= 'd0; 6505: data <= 'd2; 6506: data <= 'd1; 6507: data <= 'd1; 6508: data <= 'd1; 6509: data <= 'd3; 6510: data <= 'd6; 6511: data <= 'd6; 6512: data <= 'd6; 6513: data <= 'd6; 6514: data <= 'd6; 6515: data <= 'd3; 6516: data <= 'd1; 6517: data <= 'd1; 6518: data <= 'd2; 6519: data <= 'd0; 6520: data <= 'd0; 6521: data <= 'd0; 6522: data <= 'd0; 6523: data <= 'd0; 6524: data <= 'd0; 6525: data <= 'd0; 6526: data <= 'd0; 6527: data <= 'd0; 6528: data <= 'd0; 6529: data <= 'd0; 6530: data <= 'd0; 6531: data <= 'd0; 6532: data <= 'd0; 6533: data <= 'd0; 6534: data <= 'd0; 6535: data <= 'd0; 6536: data <= 'd0; 6537: data <= 'd2; 6538: data <= 'd1; 6539: data <= 'd1; 6540: data <= 'd5; 6541: data <= 'd5; 6542: data <= 'd5; 6543: data <= 'd1; 6544: data <= 'd1; 6545: data <= 'd1; 6546: data <= 'd1; 6547: data <= 'd1; 6548: data <= 'd5; 6549: data <= 'd5; 6550: data <= 'd2; 6551: data <= 'd0; 6552: data <= 'd0; 6553: data <= 'd0; 6554: data <= 'd0; 6555: data <= 'd0; 6556: data <= 'd0; 6557: data <= 'd0; 6558: data <= 'd0; 6559: data <= 'd0; 6560: data <= 'd0; 6561: data <= 'd0; 6562: data <= 'd0; 6563: data <= 'd0; 6564: data <= 'd0; 6565: data <= 'd0; 6566: data <= 'd0; 6567: data <= 'd0; 6568: data <= 'd2; 6569: data <= 'd1; 6570: data <= 'd5; 6571: data <= 'd5; 6572: data <= 'd3; 6573: data <= 'd6; 6574: data <= 'd6; 6575: data <= 'd6; 6576: data <= 'd6; 6577: data <= 'd6; 6578: data <= 'd6; 6579: data <= 'd6; 6580: data <= 'd6; 6581: data <= 'd3; 6582: data <= 'd5; 6583: data <= 'd2; 6584: data <= 'd0; 6585: data <= 'd0; 6586: data <= 'd0; 6587: data <= 'd0; 6588: data <= 'd0; 6589: data <= 'd0; 6590: data <= 'd0; 6591: data <= 'd0; 6592: data <= 'd0; 6593: data <= 'd0; 6594: data <= 'd0; 6595: data <= 'd0; 6596: data <= 'd0; 6597: data <= 'd0; 6598: data <= 'd0; 6599: data <= 'd0; 6600: data <= 'd2; 6601: data <= 'd5; 6602: data <= 'd3; 6603: data <= 'd6; 6604: data <= 'd3; 6605: data <= 'd1; 6606: data <= 'd1; 6607: data <= 'd1; 6608: data <= 'd1; 6609: data <= 'd1; 6610: data <= 'd1; 6611: data <= 'd1; 6612: data <= 'd1; 6613: data <= 'd1; 6614: data <= 'd3; 6615: data <= 'd2; 6616: data <= 'd0; 6617: data <= 'd0; 6618: data <= 'd0; 6619: data <= 'd0; 6620: data <= 'd0; 6621: data <= 'd0; 6622: data <= 'd0; 6623: data <= 'd0; 6624: data <= 'd0; 6625: data <= 'd0; 6626: data <= 'd0; 6627: data <= 'd0; 6628: data <= 'd0; 6629: data <= 'd0; 6630: data <= 'd0; 6631: data <= 'd0; 6632: data <= 'd2; 6633: data <= 'd5; 6634: data <= 'd3; 6635: data <= 'd1; 6636: data <= 'd1; 6637: data <= 'd1; 6638: data <= 'd5; 6639: data <= 'd5; 6640: data <= 'd5; 6641: data <= 'd5; 6642: data <= 'd5; 6643: data <= 'd5; 6644: data <= 'd5; 6645: data <= 'd1; 6646: data <= 'd1; 6647: data <= 'd2; 6648: data <= 'd0; 6649: data <= 'd0; 6650: data <= 'd0; 6651: data <= 'd0; 6652: data <= 'd0; 6653: data <= 'd0; 6654: data <= 'd0; 6655: data <= 'd0; 6656: data <= 'd0; 6657: data <= 'd0; 6658: data <= 'd0; 6659: data <= 'd0; 6660: data <= 'd0; 6661: data <= 'd0; 6662: data <= 'd2; 6663: data <= 'd2; 6664: data <= 'd2; 6665: data <= 'd6; 6666: data <= 'd1; 6667: data <= 'd5; 6668: data <= 'd2; 6669: data <= 'd2; 6670: data <= 'd2; 6671: data <= 'd2; 6672: data <= 'd2; 6673: data <= 'd2; 6674: data <= 'd2; 6675: data <= 'd2; 6676: data <= 'd2; 6677: data <= 'd2; 6678: data <= 'd5; 6679: data <= 'd2; 6680: data <= 'd0; 6681: data <= 'd0; 6682: data <= 'd0; 6683: data <= 'd0; 6684: data <= 'd0; 6685: data <= 'd0; 6686: data <= 'd0; 6687: data <= 'd0; 6688: data <= 'd0; 6689: data <= 'd0; 6690: data <= 'd0; 6691: data <= 'd0; 6692: data <= 'd0; 6693: data <= 'd0; 6694: data <= 'd2; 6695: data <= 'd1; 6696: data <= 'd2; 6697: data <= 'd1; 6698: data <= 'd5; 6699: data <= 'd2; 6700: data <= 'd8; 6701: data <= 'd8; 6702: data <= 'd8; 6703: data <= 'd8; 6704: data <= 'd8; 6705: data <= 'd9; 6706: data <= 'd9; 6707: data <= 'd8; 6708: data <= 'd8; 6709: data <= 'd8; 6710: data <= 'd2; 6711: data <= 'd2; 6712: data <= 'd0; 6713: data <= 'd0; 6714: data <= 'd0; 6715: data <= 'd0; 6716: data <= 'd0; 6717: data <= 'd0; 6718: data <= 'd0; 6719: data <= 'd0; 6720: data <= 'd0; 6721: data <= 'd0; 6722: data <= 'd0; 6723: data <= 'd0; 6724: data <= 'd0; 6725: data <= 'd0; 6726: data <= 'd2; 6727: data <= 'd5; 6728: data <= 'd2; 6729: data <= 'd1; 6730: data <= 'd2; 6731: data <= 'd8; 6732: data <= 'd8; 6733: data <= 'd9; 6734: data <= 'd9; 6735: data <= 'd2; 6736: data <= 'd9; 6737: data <= 'd11; 6738: data <= 'd11; 6739: data <= 'd10; 6740: data <= 'd2; 6741: data <= 'd9; 6742: data <= 'd2; 6743: data <= 'd2; 6744: data <= 'd0; 6745: data <= 'd0; 6746: data <= 'd0; 6747: data <= 'd0; 6748: data <= 'd0; 6749: data <= 'd0; 6750: data <= 'd0; 6751: data <= 'd0; 6752: data <= 'd0; 6753: data <= 'd0; 6754: data <= 'd0; 6755: data <= 'd0; 6756: data <= 'd0; 6757: data <= 'd0; 6758: data <= 'd0; 6759: data <= 'd2; 6760: data <= 'd5; 6761: data <= 'd2; 6762: data <= 'd9; 6763: data <= 'd10; 6764: data <= 'd9; 6765: data <= 'd9; 6766: data <= 'd10; 6767: data <= 'd11; 6768: data <= 'd10; 6769: data <= 'd11; 6770: data <= 'd11; 6771: data <= 'd10; 6772: data <= 'd11; 6773: data <= 'd10; 6774: data <= 'd9; 6775: data <= 'd2; 6776: data <= 'd0; 6777: data <= 'd0; 6778: data <= 'd0; 6779: data <= 'd0; 6780: data <= 'd0; 6781: data <= 'd0; 6782: data <= 'd0; 6783: data <= 'd0; 6784: data <= 'd0; 6785: data <= 'd0; 6786: data <= 'd0; 6787: data <= 'd0; 6788: data <= 'd0; 6789: data <= 'd0; 6790: data <= 'd0; 6791: data <= 'd0; 6792: data <= 'd2; 6793: data <= 'd2; 6794: data <= 'd2; 6795: data <= 'd8; 6796: data <= 'd9; 6797: data <= 'd9; 6798: data <= 'd10; 6799: data <= 'd10; 6800: data <= 'd10; 6801: data <= 'd8; 6802: data <= 'd8; 6803: data <= 'd10; 6804: data <= 'd10; 6805: data <= 'd9; 6806: data <= 'd2; 6807: data <= 'd0; 6808: data <= 'd0; 6809: data <= 'd0; 6810: data <= 'd0; 6811: data <= 'd0; 6812: data <= 'd0; 6813: data <= 'd0; 6814: data <= 'd0; 6815: data <= 'd0; 6816: data <= 'd0; 6817: data <= 'd0; 6818: data <= 'd0; 6819: data <= 'd0; 6820: data <= 'd0; 6821: data <= 'd0; 6822: data <= 'd0; 6823: data <= 'd0; 6824: data <= 'd0; 6825: data <= 'd0; 6826: data <= 'd2; 6827: data <= 'd8; 6828: data <= 'd8; 6829: data <= 'd9; 6830: data <= 'd9; 6831: data <= 'd10; 6832: data <= 'd10; 6833: data <= 'd9; 6834: data <= 'd9; 6835: data <= 'd10; 6836: data <= 'd10; 6837: data <= 'd9; 6838: data <= 'd2; 6839: data <= 'd0; 6840: data <= 'd0; 6841: data <= 'd0; 6842: data <= 'd0; 6843: data <= 'd0; 6844: data <= 'd0; 6845: data <= 'd0; 6846: data <= 'd0; 6847: data <= 'd0; 6848: data <= 'd0; 6849: data <= 'd0; 6850: data <= 'd0; 6851: data <= 'd0; 6852: data <= 'd0; 6853: data <= 'd0; 6854: data <= 'd0; 6855: data <= 'd0; 6856: data <= 'd0; 6857: data <= 'd0; 6858: data <= 'd2; 6859: data <= 'd2; 6860: data <= 'd5; 6861: data <= 'd5; 6862: data <= 'd8; 6863: data <= 'd9; 6864: data <= 'd9; 6865: data <= 'd9; 6866: data <= 'd9; 6867: data <= 'd9; 6868: data <= 'd9; 6869: data <= 'd5; 6870: data <= 'd2; 6871: data <= 'd0; 6872: data <= 'd0; 6873: data <= 'd0; 6874: data <= 'd0; 6875: data <= 'd0; 6876: data <= 'd0; 6877: data <= 'd0; 6878: data <= 'd0; 6879: data <= 'd0; 6880: data <= 'd0; 6881: data <= 'd0; 6882: data <= 'd0; 6883: data <= 'd0; 6884: data <= 'd0; 6885: data <= 'd0; 6886: data <= 'd0; 6887: data <= 'd0; 6888: data <= 'd0; 6889: data <= 'd2; 6890: data <= 'd7; 6891: data <= 'd1; 6892: data <= 'd1; 6893: data <= 'd1; 6894: data <= 'd3; 6895: data <= 'd3; 6896: data <= 'd3; 6897: data <= 'd5; 6898: data <= 'd5; 6899: data <= 'd3; 6900: data <= 'd3; 6901: data <= 'd1; 6902: data <= 'd2; 6903: data <= 'd0; 6904: data <= 'd0; 6905: data <= 'd0; 6906: data <= 'd0; 6907: data <= 'd0; 6908: data <= 'd0; 6909: data <= 'd0; 6910: data <= 'd0; 6911: data <= 'd0; 6912: data <= 'd0; 6913: data <= 'd0; 6914: data <= 'd0; 6915: data <= 'd0; 6916: data <= 'd0; 6917: data <= 'd0; 6918: data <= 'd0; 6919: data <= 'd0; 6920: data <= 'd0; 6921: data <= 'd2; 6922: data <= 'd7; 6923: data <= 'd7; 6924: data <= 'd1; 6925: data <= 'd1; 6926: data <= 'd3; 6927: data <= 'd3; 6928: data <= 'd3; 6929: data <= 'd1; 6930: data <= 'd1; 6931: data <= 'd3; 6932: data <= 'd3; 6933: data <= 'd1; 6934: data <= 'd2; 6935: data <= 'd0; 6936: data <= 'd0; 6937: data <= 'd0; 6938: data <= 'd0; 6939: data <= 'd0; 6940: data <= 'd0; 6941: data <= 'd0; 6942: data <= 'd0; 6943: data <= 'd0; 6944: data <= 'd0; 6945: data <= 'd0; 6946: data <= 'd0; 6947: data <= 'd0; 6948: data <= 'd0; 6949: data <= 'd0; 6950: data <= 'd0; 6951: data <= 'd0; 6952: data <= 'd0; 6953: data <= 'd2; 6954: data <= 'd9; 6955: data <= 'd9; 6956: data <= 'd5; 6957: data <= 'd1; 6958: data <= 'd1; 6959: data <= 'd3; 6960: data <= 'd3; 6961: data <= 'd1; 6962: data <= 'd1; 6963: data <= 'd3; 6964: data <= 'd1; 6965: data <= 'd1; 6966: data <= 'd8; 6967: data <= 'd2; 6968: data <= 'd0; 6969: data <= 'd0; 6970: data <= 'd0; 6971: data <= 'd0; 6972: data <= 'd0; 6973: data <= 'd0; 6974: data <= 'd0; 6975: data <= 'd0; 6976: data <= 'd0; 6977: data <= 'd0; 6978: data <= 'd0; 6979: data <= 'd0; 6980: data <= 'd0; 6981: data <= 'd0; 6982: data <= 'd0; 6983: data <= 'd0; 6984: data <= 'd0; 6985: data <= 'd2; 6986: data <= 'd9; 6987: data <= 'd9; 6988: data <= 'd2; 6989: data <= 'd2; 6990: data <= 'd2; 6991: data <= 'd2; 6992: data <= 'd5; 6993: data <= 'd5; 6994: data <= 'd5; 6995: data <= 'd2; 6996: data <= 'd2; 6997: data <= 'd2; 6998: data <= 'd8; 6999: data <= 'd2; 7000: data <= 'd0; 7001: data <= 'd0; 7002: data <= 'd0; 7003: data <= 'd0; 7004: data <= 'd0; 7005: data <= 'd0; 7006: data <= 'd0; 7007: data <= 'd0; 7008: data <= 'd0; 7009: data <= 'd0; 7010: data <= 'd0; 7011: data <= 'd0; 7012: data <= 'd0; 7013: data <= 'd0; 7014: data <= 'd0; 7015: data <= 'd0; 7016: data <= 'd0; 7017: data <= 'd0; 7018: data <= 'd2; 7019: data <= 'd2; 7020: data <= 'd1; 7021: data <= 'd1; 7022: data <= 'd3; 7023: data <= 'd3; 7024: data <= 'd3; 7025: data <= 'd1; 7026: data <= 'd3; 7027: data <= 'd3; 7028: data <= 'd3; 7029: data <= 'd2; 7030: data <= 'd2; 7031: data <= 'd0; 7032: data <= 'd0; 7033: data <= 'd0; 7034: data <= 'd0; 7035: data <= 'd0; 7036: data <= 'd0; 7037: data <= 'd0; 7038: data <= 'd0; 7039: data <= 'd0; 7040: data <= 'd0; 7041: data <= 'd0; 7042: data <= 'd0; 7043: data <= 'd0; 7044: data <= 'd0; 7045: data <= 'd0; 7046: data <= 'd0; 7047: data <= 'd0; 7048: data <= 'd0; 7049: data <= 'd0; 7050: data <= 'd0; 7051: data <= 'd2; 7052: data <= 'd4; 7053: data <= 'd7; 7054: data <= 'd7; 7055: data <= 'd2; 7056: data <= 'd2; 7057: data <= 'd2; 7058: data <= 'd5; 7059: data <= 'd5; 7060: data <= 'd4; 7061: data <= 'd2; 7062: data <= 'd0; 7063: data <= 'd0; 7064: data <= 'd0; 7065: data <= 'd0; 7066: data <= 'd0; 7067: data <= 'd0; 7068: data <= 'd0; 7069: data <= 'd0; 7070: data <= 'd0; 7071: data <= 'd0; 7072: data <= 'd0; 7073: data <= 'd0; 7074: data <= 'd0; 7075: data <= 'd0; 7076: data <= 'd0; 7077: data <= 'd0; 7078: data <= 'd0; 7079: data <= 'd0; 7080: data <= 'd0; 7081: data <= 'd0; 7082: data <= 'd0; 7083: data <= 'd0; 7084: data <= 'd2; 7085: data <= 'd4; 7086: data <= 'd7; 7087: data <= 'd2; 7088: data <= 'd0; 7089: data <= 'd0; 7090: data <= 'd2; 7091: data <= 'd4; 7092: data <= 'd4; 7093: data <= 'd2; 7094: data <= 'd0; 7095: data <= 'd0; 7096: data <= 'd0; 7097: data <= 'd0; 7098: data <= 'd0; 7099: data <= 'd0; 7100: data <= 'd0; 7101: data <= 'd0; 7102: data <= 'd0; 7103: data <= 'd0; 7104: data <= 'd0; 7105: data <= 'd0; 7106: data <= 'd0; 7107: data <= 'd0; 7108: data <= 'd0; 7109: data <= 'd0; 7110: data <= 'd0; 7111: data <= 'd0; 7112: data <= 'd0; 7113: data <= 'd0; 7114: data <= 'd0; 7115: data <= 'd0; 7116: data <= 'd2; 7117: data <= 'd2; 7118: data <= 'd2; 7119: data <= 'd0; 7120: data <= 'd0; 7121: data <= 'd0; 7122: data <= 'd0; 7123: data <= 'd2; 7124: data <= 'd2; 7125: data <= 'd2; 7126: data <= 'd0; 7127: data <= 'd0; 7128: data <= 'd0; 7129: data <= 'd0; 7130: data <= 'd0; 7131: data <= 'd0; 7132: data <= 'd0; 7133: data <= 'd0; 7134: data <= 'd0; 7135: data <= 'd0; 7136: data <= 'd0; 7137: data <= 'd0; 7138: data <= 'd0; 7139: data <= 'd0; 7140: data <= 'd0; 7141: data <= 'd0; 7142: data <= 'd0; 7143: data <= 'd0; 7144: data <= 'd0; 7145: data <= 'd0; 7146: data <= 'd0; 7147: data <= 'd0; 7148: data <= 'd0; 7149: data <= 'd0; 7150: data <= 'd0; 7151: data <= 'd0; 7152: data <= 'd0; 7153: data <= 'd0; 7154: data <= 'd0; 7155: data <= 'd0; 7156: data <= 'd0; 7157: data <= 'd0; 7158: data <= 'd0; 7159: data <= 'd0; 7160: data <= 'd0; 7161: data <= 'd0; 7162: data <= 'd0; 7163: data <= 'd0; 7164: data <= 'd0; 7165: data <= 'd0; 7166: data <= 'd0; 7167: data <= 'd0; 7168: data <= 'd0; 7169: data <= 'd0; 7170: data <= 'd0; 7171: data <= 'd0; 7172: data <= 'd0; 7173: data <= 'd0; 7174: data <= 'd0; 7175: data <= 'd0; 7176: data <= 'd0; 7177: data <= 'd0; 7178: data <= 'd0; 7179: data <= 'd0; 7180: data <= 'd0; 7181: data <= 'd0; 7182: data <= 'd0; 7183: data <= 'd0; 7184: data <= 'd0; 7185: data <= 'd0; 7186: data <= 'd0; 7187: data <= 'd0; 7188: data <= 'd0; 7189: data <= 'd0; 7190: data <= 'd0; 7191: data <= 'd0; 7192: data <= 'd0; 7193: data <= 'd0; 7194: data <= 'd0; 7195: data <= 'd0; 7196: data <= 'd0; 7197: data <= 'd0; 7198: data <= 'd0; 7199: data <= 'd0; 7200: data <= 'd0; 7201: data <= 'd0; 7202: data <= 'd0; 7203: data <= 'd0; 7204: data <= 'd0; 7205: data <= 'd0; 7206: data <= 'd0; 7207: data <= 'd0; 7208: data <= 'd0; 7209: data <= 'd0; 7210: data <= 'd0; 7211: data <= 'd0; 7212: data <= 'd0; 7213: data <= 'd0; 7214: data <= 'd0; 7215: data <= 'd0; 7216: data <= 'd0; 7217: data <= 'd0; 7218: data <= 'd0; 7219: data <= 'd0; 7220: data <= 'd0; 7221: data <= 'd0; 7222: data <= 'd0; 7223: data <= 'd0; 7224: data <= 'd0; 7225: data <= 'd0; 7226: data <= 'd0; 7227: data <= 'd0; 7228: data <= 'd0; 7229: data <= 'd0; 7230: data <= 'd0; 7231: data <= 'd0; 7232: data <= 'd0; 7233: data <= 'd0; 7234: data <= 'd0; 7235: data <= 'd0; 7236: data <= 'd0; 7237: data <= 'd0; 7238: data <= 'd0; 7239: data <= 'd0; 7240: data <= 'd0; 7241: data <= 'd0; 7242: data <= 'd0; 7243: data <= 'd0; 7244: data <= 'd0; 7245: data <= 'd0; 7246: data <= 'd0; 7247: data <= 'd0; 7248: data <= 'd0; 7249: data <= 'd0; 7250: data <= 'd0; 7251: data <= 'd0; 7252: data <= 'd0; 7253: data <= 'd0; 7254: data <= 'd0; 7255: data <= 'd0; 7256: data <= 'd0; 7257: data <= 'd0; 7258: data <= 'd0; 7259: data <= 'd0; 7260: data <= 'd0; 7261: data <= 'd0; 7262: data <= 'd0; 7263: data <= 'd0; 7264: data <= 'd0; 7265: data <= 'd0; 7266: data <= 'd0; 7267: data <= 'd0; 7268: data <= 'd0; 7269: data <= 'd0; 7270: data <= 'd0; 7271: data <= 'd0; 7272: data <= 'd0; 7273: data <= 'd0; 7274: data <= 'd0; 7275: data <= 'd0; 7276: data <= 'd0; 7277: data <= 'd0; 7278: data <= 'd0; 7279: data <= 'd0; 7280: data <= 'd0; 7281: data <= 'd0; 7282: data <= 'd0; 7283: data <= 'd0; 7284: data <= 'd0; 7285: data <= 'd0; 7286: data <= 'd0; 7287: data <= 'd0; 7288: data <= 'd0; 7289: data <= 'd0; 7290: data <= 'd0; 7291: data <= 'd0; 7292: data <= 'd0; 7293: data <= 'd0; 7294: data <= 'd0; 7295: data <= 'd0; 7296: data <= 'd0; 7297: data <= 'd0; 7298: data <= 'd0; 7299: data <= 'd0; 7300: data <= 'd0; 7301: data <= 'd0; 7302: data <= 'd0; 7303: data <= 'd0; 7304: data <= 'd0; 7305: data <= 'd0; 7306: data <= 'd0; 7307: data <= 'd0; 7308: data <= 'd0; 7309: data <= 'd0; 7310: data <= 'd0; 7311: data <= 'd0; 7312: data <= 'd0; 7313: data <= 'd0; 7314: data <= 'd0; 7315: data <= 'd0; 7316: data <= 'd0; 7317: data <= 'd0; 7318: data <= 'd0; 7319: data <= 'd0; 7320: data <= 'd0; 7321: data <= 'd0; 7322: data <= 'd0; 7323: data <= 'd0; 7324: data <= 'd0; 7325: data <= 'd0; 7326: data <= 'd0; 7327: data <= 'd0; 7328: data <= 'd0; 7329: data <= 'd0; 7330: data <= 'd0; 7331: data <= 'd0; 7332: data <= 'd0; 7333: data <= 'd0; 7334: data <= 'd0; 7335: data <= 'd0; 7336: data <= 'd0; 7337: data <= 'd0; 7338: data <= 'd0; 7339: data <= 'd0; 7340: data <= 'd0; 7341: data <= 'd0; 7342: data <= 'd0; 7343: data <= 'd0; 7344: data <= 'd0; 7345: data <= 'd0; 7346: data <= 'd0; 7347: data <= 'd0; 7348: data <= 'd0; 7349: data <= 'd0; 7350: data <= 'd0; 7351: data <= 'd0; 7352: data <= 'd0; 7353: data <= 'd0; 7354: data <= 'd0; 7355: data <= 'd0; 7356: data <= 'd0; 7357: data <= 'd0; 7358: data <= 'd0; 7359: data <= 'd0; 7360: data <= 'd0; 7361: data <= 'd0; 7362: data <= 'd0; 7363: data <= 'd0; 7364: data <= 'd0; 7365: data <= 'd0; 7366: data <= 'd0; 7367: data <= 'd0; 7368: data <= 'd0; 7369: data <= 'd0; 7370: data <= 'd0; 7371: data <= 'd0; 7372: data <= 'd0; 7373: data <= 'd0; 7374: data <= 'd0; 7375: data <= 'd0; 7376: data <= 'd0; 7377: data <= 'd0; 7378: data <= 'd0; 7379: data <= 'd0; 7380: data <= 'd0; 7381: data <= 'd0; 7382: data <= 'd0; 7383: data <= 'd0; 7384: data <= 'd0; 7385: data <= 'd0; 7386: data <= 'd0; 7387: data <= 'd0; 7388: data <= 'd0; 7389: data <= 'd0; 7390: data <= 'd0; 7391: data <= 'd0; 7392: data <= 'd0; 7393: data <= 'd0; 7394: data <= 'd0; 7395: data <= 'd0; 7396: data <= 'd0; 7397: data <= 'd0; 7398: data <= 'd0; 7399: data <= 'd0; 7400: data <= 'd0; 7401: data <= 'd0; 7402: data <= 'd0; 7403: data <= 'd0; 7404: data <= 'd0; 7405: data <= 'd0; 7406: data <= 'd0; 7407: data <= 'd0; 7408: data <= 'd0; 7409: data <= 'd0; 7410: data <= 'd0; 7411: data <= 'd0; 7412: data <= 'd0; 7413: data <= 'd0; 7414: data <= 'd0; 7415: data <= 'd0; 7416: data <= 'd0; 7417: data <= 'd0; 7418: data <= 'd0; 7419: data <= 'd0; 7420: data <= 'd0; 7421: data <= 'd0; 7422: data <= 'd0; 7423: data <= 'd0; 7424: data <= 'd0; 7425: data <= 'd0; 7426: data <= 'd0; 7427: data <= 'd0; 7428: data <= 'd0; 7429: data <= 'd0; 7430: data <= 'd0; 7431: data <= 'd0; 7432: data <= 'd0; 7433: data <= 'd0; 7434: data <= 'd0; 7435: data <= 'd0; 7436: data <= 'd0; 7437: data <= 'd0; 7438: data <= 'd0; 7439: data <= 'd0; 7440: data <= 'd0; 7441: data <= 'd0; 7442: data <= 'd0; 7443: data <= 'd0; 7444: data <= 'd0; 7445: data <= 'd0; 7446: data <= 'd0; 7447: data <= 'd0; 7448: data <= 'd0; 7449: data <= 'd0; 7450: data <= 'd0; 7451: data <= 'd0; 7452: data <= 'd0; 7453: data <= 'd0; 7454: data <= 'd0; 7455: data <= 'd0; 7456: data <= 'd0; 7457: data <= 'd0; 7458: data <= 'd0; 7459: data <= 'd0; 7460: data <= 'd0; 7461: data <= 'd0; 7462: data <= 'd0; 7463: data <= 'd0; 7464: data <= 'd0; 7465: data <= 'd0; 7466: data <= 'd0; 7467: data <= 'd0; 7468: data <= 'd0; 7469: data <= 'd0; 7470: data <= 'd0; 7471: data <= 'd0; 7472: data <= 'd0; 7473: data <= 'd0; 7474: data <= 'd0; 7475: data <= 'd0; 7476: data <= 'd0; 7477: data <= 'd0; 7478: data <= 'd0; 7479: data <= 'd0; 7480: data <= 'd0; 7481: data <= 'd0; 7482: data <= 'd0; 7483: data <= 'd0; 7484: data <= 'd0; 7485: data <= 'd0; 7486: data <= 'd0; 7487: data <= 'd0; 7488: data <= 'd0; 7489: data <= 'd0; 7490: data <= 'd0; 7491: data <= 'd0; 7492: data <= 'd0; 7493: data <= 'd0; 7494: data <= 'd0; 7495: data <= 'd0; 7496: data <= 'd0; 7497: data <= 'd0; 7498: data <= 'd0; 7499: data <= 'd0; 7500: data <= 'd0; 7501: data <= 'd2; 7502: data <= 'd2; 7503: data <= 'd2; 7504: data <= 'd2; 7505: data <= 'd2; 7506: data <= 'd2; 7507: data <= 'd0; 7508: data <= 'd0; 7509: data <= 'd0; 7510: data <= 'd0; 7511: data <= 'd0; 7512: data <= 'd0; 7513: data <= 'd0; 7514: data <= 'd0; 7515: data <= 'd0; 7516: data <= 'd0; 7517: data <= 'd0; 7518: data <= 'd0; 7519: data <= 'd0; 7520: data <= 'd0; 7521: data <= 'd0; 7522: data <= 'd0; 7523: data <= 'd0; 7524: data <= 'd0; 7525: data <= 'd0; 7526: data <= 'd0; 7527: data <= 'd0; 7528: data <= 'd0; 7529: data <= 'd0; 7530: data <= 'd0; 7531: data <= 'd2; 7532: data <= 'd2; 7533: data <= 'd6; 7534: data <= 'd6; 7535: data <= 'd6; 7536: data <= 'd6; 7537: data <= 'd6; 7538: data <= 'd6; 7539: data <= 'd2; 7540: data <= 'd2; 7541: data <= 'd0; 7542: data <= 'd0; 7543: data <= 'd0; 7544: data <= 'd0; 7545: data <= 'd0; 7546: data <= 'd0; 7547: data <= 'd0; 7548: data <= 'd0; 7549: data <= 'd0; 7550: data <= 'd0; 7551: data <= 'd0; 7552: data <= 'd0; 7553: data <= 'd0; 7554: data <= 'd0; 7555: data <= 'd0; 7556: data <= 'd0; 7557: data <= 'd0; 7558: data <= 'd0; 7559: data <= 'd0; 7560: data <= 'd0; 7561: data <= 'd0; 7562: data <= 'd2; 7563: data <= 'd1; 7564: data <= 'd3; 7565: data <= 'd6; 7566: data <= 'd6; 7567: data <= 'd6; 7568: data <= 'd6; 7569: data <= 'd6; 7570: data <= 'd6; 7571: data <= 'd6; 7572: data <= 'd3; 7573: data <= 'd2; 7574: data <= 'd0; 7575: data <= 'd0; 7576: data <= 'd0; 7577: data <= 'd0; 7578: data <= 'd0; 7579: data <= 'd0; 7580: data <= 'd0; 7581: data <= 'd0; 7582: data <= 'd0; 7583: data <= 'd0; 7584: data <= 'd0; 7585: data <= 'd0; 7586: data <= 'd0; 7587: data <= 'd0; 7588: data <= 'd0; 7589: data <= 'd0; 7590: data <= 'd0; 7591: data <= 'd0; 7592: data <= 'd0; 7593: data <= 'd2; 7594: data <= 'd1; 7595: data <= 'd1; 7596: data <= 'd1; 7597: data <= 'd3; 7598: data <= 'd6; 7599: data <= 'd6; 7600: data <= 'd6; 7601: data <= 'd6; 7602: data <= 'd6; 7603: data <= 'd3; 7604: data <= 'd1; 7605: data <= 'd1; 7606: data <= 'd2; 7607: data <= 'd0; 7608: data <= 'd0; 7609: data <= 'd0; 7610: data <= 'd0; 7611: data <= 'd0; 7612: data <= 'd0; 7613: data <= 'd0; 7614: data <= 'd0; 7615: data <= 'd0; 7616: data <= 'd0; 7617: data <= 'd0; 7618: data <= 'd0; 7619: data <= 'd0; 7620: data <= 'd0; 7621: data <= 'd0; 7622: data <= 'd0; 7623: data <= 'd0; 7624: data <= 'd0; 7625: data <= 'd2; 7626: data <= 'd1; 7627: data <= 'd1; 7628: data <= 'd5; 7629: data <= 'd5; 7630: data <= 'd5; 7631: data <= 'd1; 7632: data <= 'd1; 7633: data <= 'd1; 7634: data <= 'd1; 7635: data <= 'd1; 7636: data <= 'd5; 7637: data <= 'd5; 7638: data <= 'd2; 7639: data <= 'd0; 7640: data <= 'd0; 7641: data <= 'd0; 7642: data <= 'd0; 7643: data <= 'd0; 7644: data <= 'd0; 7645: data <= 'd0; 7646: data <= 'd0; 7647: data <= 'd0; 7648: data <= 'd0; 7649: data <= 'd0; 7650: data <= 'd0; 7651: data <= 'd0; 7652: data <= 'd0; 7653: data <= 'd0; 7654: data <= 'd0; 7655: data <= 'd0; 7656: data <= 'd2; 7657: data <= 'd1; 7658: data <= 'd5; 7659: data <= 'd5; 7660: data <= 'd3; 7661: data <= 'd6; 7662: data <= 'd6; 7663: data <= 'd6; 7664: data <= 'd6; 7665: data <= 'd6; 7666: data <= 'd6; 7667: data <= 'd6; 7668: data <= 'd6; 7669: data <= 'd3; 7670: data <= 'd5; 7671: data <= 'd2; 7672: data <= 'd0; 7673: data <= 'd0; 7674: data <= 'd0; 7675: data <= 'd0; 7676: data <= 'd0; 7677: data <= 'd0; 7678: data <= 'd0; 7679: data <= 'd0; 7680: data <= 'd0; 7681: data <= 'd0; 7682: data <= 'd0; 7683: data <= 'd0; 7684: data <= 'd0; 7685: data <= 'd0; 7686: data <= 'd0; 7687: data <= 'd0; 7688: data <= 'd2; 7689: data <= 'd5; 7690: data <= 'd3; 7691: data <= 'd6; 7692: data <= 'd3; 7693: data <= 'd1; 7694: data <= 'd1; 7695: data <= 'd1; 7696: data <= 'd1; 7697: data <= 'd1; 7698: data <= 'd1; 7699: data <= 'd1; 7700: data <= 'd1; 7701: data <= 'd1; 7702: data <= 'd3; 7703: data <= 'd2; 7704: data <= 'd0; 7705: data <= 'd0; 7706: data <= 'd0; 7707: data <= 'd0; 7708: data <= 'd0; 7709: data <= 'd0; 7710: data <= 'd0; 7711: data <= 'd0; 7712: data <= 'd0; 7713: data <= 'd0; 7714: data <= 'd0; 7715: data <= 'd0; 7716: data <= 'd0; 7717: data <= 'd0; 7718: data <= 'd0; 7719: data <= 'd0; 7720: data <= 'd2; 7721: data <= 'd5; 7722: data <= 'd3; 7723: data <= 'd1; 7724: data <= 'd1; 7725: data <= 'd1; 7726: data <= 'd5; 7727: data <= 'd5; 7728: data <= 'd5; 7729: data <= 'd5; 7730: data <= 'd5; 7731: data <= 'd5; 7732: data <= 'd5; 7733: data <= 'd1; 7734: data <= 'd1; 7735: data <= 'd2; 7736: data <= 'd0; 7737: data <= 'd0; 7738: data <= 'd0; 7739: data <= 'd0; 7740: data <= 'd0; 7741: data <= 'd0; 7742: data <= 'd0; 7743: data <= 'd0; 7744: data <= 'd0; 7745: data <= 'd0; 7746: data <= 'd0; 7747: data <= 'd0; 7748: data <= 'd0; 7749: data <= 'd0; 7750: data <= 'd0; 7751: data <= 'd0; 7752: data <= 'd2; 7753: data <= 'd6; 7754: data <= 'd1; 7755: data <= 'd5; 7756: data <= 'd2; 7757: data <= 'd2; 7758: data <= 'd2; 7759: data <= 'd2; 7760: data <= 'd2; 7761: data <= 'd2; 7762: data <= 'd2; 7763: data <= 'd2; 7764: data <= 'd2; 7765: data <= 'd2; 7766: data <= 'd5; 7767: data <= 'd2; 7768: data <= 'd0; 7769: data <= 'd0; 7770: data <= 'd0; 7771: data <= 'd0; 7772: data <= 'd0; 7773: data <= 'd0; 7774: data <= 'd0; 7775: data <= 'd0; 7776: data <= 'd0; 7777: data <= 'd0; 7778: data <= 'd0; 7779: data <= 'd0; 7780: data <= 'd0; 7781: data <= 'd0; 7782: data <= 'd2; 7783: data <= 'd2; 7784: data <= 'd2; 7785: data <= 'd1; 7786: data <= 'd5; 7787: data <= 'd2; 7788: data <= 'd8; 7789: data <= 'd8; 7790: data <= 'd8; 7791: data <= 'd8; 7792: data <= 'd8; 7793: data <= 'd9; 7794: data <= 'd9; 7795: data <= 'd8; 7796: data <= 'd8; 7797: data <= 'd8; 7798: data <= 'd2; 7799: data <= 'd2; 7800: data <= 'd0; 7801: data <= 'd0; 7802: data <= 'd0; 7803: data <= 'd0; 7804: data <= 'd0; 7805: data <= 'd0; 7806: data <= 'd0; 7807: data <= 'd0; 7808: data <= 'd0; 7809: data <= 'd0; 7810: data <= 'd0; 7811: data <= 'd0; 7812: data <= 'd0; 7813: data <= 'd0; 7814: data <= 'd2; 7815: data <= 'd1; 7816: data <= 'd2; 7817: data <= 'd1; 7818: data <= 'd2; 7819: data <= 'd8; 7820: data <= 'd8; 7821: data <= 'd9; 7822: data <= 'd9; 7823: data <= 'd2; 7824: data <= 'd9; 7825: data <= 'd11; 7826: data <= 'd11; 7827: data <= 'd10; 7828: data <= 'd2; 7829: data <= 'd9; 7830: data <= 'd2; 7831: data <= 'd2; 7832: data <= 'd0; 7833: data <= 'd0; 7834: data <= 'd0; 7835: data <= 'd0; 7836: data <= 'd0; 7837: data <= 'd0; 7838: data <= 'd0; 7839: data <= 'd0; 7840: data <= 'd0; 7841: data <= 'd0; 7842: data <= 'd0; 7843: data <= 'd0; 7844: data <= 'd0; 7845: data <= 'd0; 7846: data <= 'd2; 7847: data <= 'd5; 7848: data <= 'd1; 7849: data <= 'd2; 7850: data <= 'd9; 7851: data <= 'd10; 7852: data <= 'd9; 7853: data <= 'd9; 7854: data <= 'd10; 7855: data <= 'd11; 7856: data <= 'd10; 7857: data <= 'd11; 7858: data <= 'd11; 7859: data <= 'd10; 7860: data <= 'd11; 7861: data <= 'd10; 7862: data <= 'd9; 7863: data <= 'd2; 7864: data <= 'd0; 7865: data <= 'd0; 7866: data <= 'd0; 7867: data <= 'd0; 7868: data <= 'd0; 7869: data <= 'd0; 7870: data <= 'd0; 7871: data <= 'd0; 7872: data <= 'd0; 7873: data <= 'd0; 7874: data <= 'd0; 7875: data <= 'd0; 7876: data <= 'd0; 7877: data <= 'd0; 7878: data <= 'd0; 7879: data <= 'd2; 7880: data <= 'd5; 7881: data <= 'd5; 7882: data <= 'd2; 7883: data <= 'd8; 7884: data <= 'd9; 7885: data <= 'd9; 7886: data <= 'd10; 7887: data <= 'd10; 7888: data <= 'd10; 7889: data <= 'd8; 7890: data <= 'd8; 7891: data <= 'd10; 7892: data <= 'd10; 7893: data <= 'd9; 7894: data <= 'd2; 7895: data <= 'd0; 7896: data <= 'd0; 7897: data <= 'd0; 7898: data <= 'd0; 7899: data <= 'd0; 7900: data <= 'd0; 7901: data <= 'd0; 7902: data <= 'd0; 7903: data <= 'd0; 7904: data <= 'd0; 7905: data <= 'd0; 7906: data <= 'd0; 7907: data <= 'd0; 7908: data <= 'd0; 7909: data <= 'd0; 7910: data <= 'd0; 7911: data <= 'd0; 7912: data <= 'd2; 7913: data <= 'd2; 7914: data <= 'd2; 7915: data <= 'd8; 7916: data <= 'd8; 7917: data <= 'd9; 7918: data <= 'd9; 7919: data <= 'd10; 7920: data <= 'd10; 7921: data <= 'd9; 7922: data <= 'd9; 7923: data <= 'd10; 7924: data <= 'd10; 7925: data <= 'd9; 7926: data <= 'd2; 7927: data <= 'd0; 7928: data <= 'd0; 7929: data <= 'd0; 7930: data <= 'd0; 7931: data <= 'd0; 7932: data <= 'd0; 7933: data <= 'd0; 7934: data <= 'd0; 7935: data <= 'd0; 7936: data <= 'd0; 7937: data <= 'd0; 7938: data <= 'd0; 7939: data <= 'd0; 7940: data <= 'd0; 7941: data <= 'd0; 7942: data <= 'd0; 7943: data <= 'd0; 7944: data <= 'd0; 7945: data <= 'd0; 7946: data <= 'd2; 7947: data <= 'd2; 7948: data <= 'd5; 7949: data <= 'd5; 7950: data <= 'd8; 7951: data <= 'd9; 7952: data <= 'd9; 7953: data <= 'd9; 7954: data <= 'd9; 7955: data <= 'd9; 7956: data <= 'd9; 7957: data <= 'd5; 7958: data <= 'd2; 7959: data <= 'd0; 7960: data <= 'd0; 7961: data <= 'd0; 7962: data <= 'd0; 7963: data <= 'd0; 7964: data <= 'd0; 7965: data <= 'd0; 7966: data <= 'd0; 7967: data <= 'd0; 7968: data <= 'd0; 7969: data <= 'd0; 7970: data <= 'd0; 7971: data <= 'd0; 7972: data <= 'd0; 7973: data <= 'd0; 7974: data <= 'd0; 7975: data <= 'd0; 7976: data <= 'd0; 7977: data <= 'd2; 7978: data <= 'd7; 7979: data <= 'd1; 7980: data <= 'd1; 7981: data <= 'd1; 7982: data <= 'd3; 7983: data <= 'd3; 7984: data <= 'd3; 7985: data <= 'd5; 7986: data <= 'd5; 7987: data <= 'd3; 7988: data <= 'd3; 7989: data <= 'd1; 7990: data <= 'd2; 7991: data <= 'd0; 7992: data <= 'd0; 7993: data <= 'd0; 7994: data <= 'd0; 7995: data <= 'd0; 7996: data <= 'd0; 7997: data <= 'd0; 7998: data <= 'd0; 7999: data <= 'd0; 8000: data <= 'd0; 8001: data <= 'd0; 8002: data <= 'd0; 8003: data <= 'd0; 8004: data <= 'd0; 8005: data <= 'd0; 8006: data <= 'd0; 8007: data <= 'd0; 8008: data <= 'd0; 8009: data <= 'd2; 8010: data <= 'd7; 8011: data <= 'd7; 8012: data <= 'd5; 8013: data <= 'd1; 8014: data <= 'd3; 8015: data <= 'd3; 8016: data <= 'd3; 8017: data <= 'd1; 8018: data <= 'd1; 8019: data <= 'd3; 8020: data <= 'd3; 8021: data <= 'd1; 8022: data <= 'd2; 8023: data <= 'd2; 8024: data <= 'd0; 8025: data <= 'd0; 8026: data <= 'd0; 8027: data <= 'd0; 8028: data <= 'd0; 8029: data <= 'd0; 8030: data <= 'd0; 8031: data <= 'd0; 8032: data <= 'd0; 8033: data <= 'd0; 8034: data <= 'd0; 8035: data <= 'd0; 8036: data <= 'd0; 8037: data <= 'd0; 8038: data <= 'd0; 8039: data <= 'd0; 8040: data <= 'd0; 8041: data <= 'd0; 8042: data <= 'd2; 8043: data <= 'd9; 8044: data <= 'd9; 8045: data <= 'd2; 8046: data <= 'd1; 8047: data <= 'd3; 8048: data <= 'd3; 8049: data <= 'd1; 8050: data <= 'd1; 8051: data <= 'd3; 8052: data <= 'd1; 8053: data <= 'd1; 8054: data <= 'd8; 8055: data <= 'd9; 8056: data <= 'd2; 8057: data <= 'd0; 8058: data <= 'd0; 8059: data <= 'd0; 8060: data <= 'd0; 8061: data <= 'd0; 8062: data <= 'd0; 8063: data <= 'd0; 8064: data <= 'd0; 8065: data <= 'd0; 8066: data <= 'd0; 8067: data <= 'd0; 8068: data <= 'd0; 8069: data <= 'd0; 8070: data <= 'd0; 8071: data <= 'd0; 8072: data <= 'd0; 8073: data <= 'd0; 8074: data <= 'd2; 8075: data <= 'd9; 8076: data <= 'd9; 8077: data <= 'd2; 8078: data <= 'd2; 8079: data <= 'd2; 8080: data <= 'd5; 8081: data <= 'd5; 8082: data <= 'd5; 8083: data <= 'd2; 8084: data <= 'd2; 8085: data <= 'd2; 8086: data <= 'd8; 8087: data <= 'd9; 8088: data <= 'd2; 8089: data <= 'd0; 8090: data <= 'd0; 8091: data <= 'd0; 8092: data <= 'd0; 8093: data <= 'd0; 8094: data <= 'd0; 8095: data <= 'd0; 8096: data <= 'd0; 8097: data <= 'd0; 8098: data <= 'd0; 8099: data <= 'd0; 8100: data <= 'd0; 8101: data <= 'd0; 8102: data <= 'd0; 8103: data <= 'd0; 8104: data <= 'd0; 8105: data <= 'd0; 8106: data <= 'd0; 8107: data <= 'd2; 8108: data <= 'd2; 8109: data <= 'd1; 8110: data <= 'd3; 8111: data <= 'd3; 8112: data <= 'd3; 8113: data <= 'd1; 8114: data <= 'd3; 8115: data <= 'd3; 8116: data <= 'd3; 8117: data <= 'd2; 8118: data <= 'd2; 8119: data <= 'd2; 8120: data <= 'd0; 8121: data <= 'd0; 8122: data <= 'd0; 8123: data <= 'd0; 8124: data <= 'd0; 8125: data <= 'd0; 8126: data <= 'd0; 8127: data <= 'd0; 8128: data <= 'd0; 8129: data <= 'd0; 8130: data <= 'd0; 8131: data <= 'd0; 8132: data <= 'd0; 8133: data <= 'd0; 8134: data <= 'd0; 8135: data <= 'd0; 8136: data <= 'd0; 8137: data <= 'd0; 8138: data <= 'd0; 8139: data <= 'd2; 8140: data <= 'd4; 8141: data <= 'd7; 8142: data <= 'd7; 8143: data <= 'd2; 8144: data <= 'd2; 8145: data <= 'd2; 8146: data <= 'd5; 8147: data <= 'd5; 8148: data <= 'd4; 8149: data <= 'd2; 8150: data <= 'd0; 8151: data <= 'd0; 8152: data <= 'd0; 8153: data <= 'd0; 8154: data <= 'd0; 8155: data <= 'd0; 8156: data <= 'd0; 8157: data <= 'd0; 8158: data <= 'd0; 8159: data <= 'd0; 8160: data <= 'd0; 8161: data <= 'd0; 8162: data <= 'd0; 8163: data <= 'd0; 8164: data <= 'd0; 8165: data <= 'd0; 8166: data <= 'd0; 8167: data <= 'd0; 8168: data <= 'd0; 8169: data <= 'd0; 8170: data <= 'd0; 8171: data <= 'd0; 8172: data <= 'd2; 8173: data <= 'd2; 8174: data <= 'd2; 8175: data <= 'd0; 8176: data <= 'd0; 8177: data <= 'd0; 8178: data <= 'd2; 8179: data <= 'd2; 8180: data <= 'd2; 8181: data <= 'd0; 8182: data <= 'd0; 8183: data <= 'd0; 8184: data <= 'd0; 8185: data <= 'd0; 8186: data <= 'd0; 8187: data <= 'd0; 8188: data <= 'd0; 8189: data <= 'd0; 8190: data <= 'd0; 8191: data <= 'd0; 8192: data <= 'd0; 8193: data <= 'd0; 8194: data <= 'd0; 8195: data <= 'd0; 8196: data <= 'd0; 8197: data <= 'd0; 8198: data <= 'd0; 8199: data <= 'd0; 8200: data <= 'd0; 8201: data <= 'd0; 8202: data <= 'd0; 8203: data <= 'd0; 8204: data <= 'd0; 8205: data <= 'd0; 8206: data <= 'd0; 8207: data <= 'd0; 8208: data <= 'd0; 8209: data <= 'd0; 8210: data <= 'd0; 8211: data <= 'd0; 8212: data <= 'd0; 8213: data <= 'd0; 8214: data <= 'd0; 8215: data <= 'd0; 8216: data <= 'd0; 8217: data <= 'd0; 8218: data <= 'd0; 8219: data <= 'd0; 8220: data <= 'd0; 8221: data <= 'd0; 8222: data <= 'd0; 8223: data <= 'd0; 8224: data <= 'd0; 8225: data <= 'd0; 8226: data <= 'd0; 8227: data <= 'd0; 8228: data <= 'd0; 8229: data <= 'd0; 8230: data <= 'd0; 8231: data <= 'd0; 8232: data <= 'd0; 8233: data <= 'd0; 8234: data <= 'd0; 8235: data <= 'd0; 8236: data <= 'd0; 8237: data <= 'd0; 8238: data <= 'd0; 8239: data <= 'd0; 8240: data <= 'd0; 8241: data <= 'd0; 8242: data <= 'd0; 8243: data <= 'd0; 8244: data <= 'd0; 8245: data <= 'd0; 8246: data <= 'd0; 8247: data <= 'd0; 8248: data <= 'd0; 8249: data <= 'd0; 8250: data <= 'd0; 8251: data <= 'd0; 8252: data <= 'd0; 8253: data <= 'd0; 8254: data <= 'd0; 8255: data <= 'd0; 8256: data <= 'd0; 8257: data <= 'd0; 8258: data <= 'd0; 8259: data <= 'd0; 8260: data <= 'd0; 8261: data <= 'd0; 8262: data <= 'd0; 8263: data <= 'd0; 8264: data <= 'd0; 8265: data <= 'd0; 8266: data <= 'd0; 8267: data <= 'd0; 8268: data <= 'd0; 8269: data <= 'd0; 8270: data <= 'd0; 8271: data <= 'd0; 8272: data <= 'd0; 8273: data <= 'd0; 8274: data <= 'd0; 8275: data <= 'd0; 8276: data <= 'd0; 8277: data <= 'd0; 8278: data <= 'd0; 8279: data <= 'd0; 8280: data <= 'd0; 8281: data <= 'd0; 8282: data <= 'd0; 8283: data <= 'd0; 8284: data <= 'd0; 8285: data <= 'd0; 8286: data <= 'd0; 8287: data <= 'd0; 8288: data <= 'd0; 8289: data <= 'd0; 8290: data <= 'd0; 8291: data <= 'd0; 8292: data <= 'd0; 8293: data <= 'd0; 8294: data <= 'd0; 8295: data <= 'd0; 8296: data <= 'd0; 8297: data <= 'd0; 8298: data <= 'd0; 8299: data <= 'd0; 8300: data <= 'd0; 8301: data <= 'd0; 8302: data <= 'd0; 8303: data <= 'd0; 8304: data <= 'd0; 8305: data <= 'd0; 8306: data <= 'd0; 8307: data <= 'd0; 8308: data <= 'd0; 8309: data <= 'd0; 8310: data <= 'd0; 8311: data <= 'd0; 8312: data <= 'd0; 8313: data <= 'd0; 8314: data <= 'd0; 8315: data <= 'd0; 8316: data <= 'd0; 8317: data <= 'd0; 8318: data <= 'd0; 8319: data <= 'd0; 8320: data <= 'd0; 8321: data <= 'd0; 8322: data <= 'd0; 8323: data <= 'd0; 8324: data <= 'd0; 8325: data <= 'd0; 8326: data <= 'd0; 8327: data <= 'd0; 8328: data <= 'd0; 8329: data <= 'd0; 8330: data <= 'd0; 8331: data <= 'd0; 8332: data <= 'd0; 8333: data <= 'd0; 8334: data <= 'd0; 8335: data <= 'd0; 8336: data <= 'd0; 8337: data <= 'd0; 8338: data <= 'd0; 8339: data <= 'd0; 8340: data <= 'd0; 8341: data <= 'd0; 8342: data <= 'd0; 8343: data <= 'd0; 8344: data <= 'd0; 8345: data <= 'd0; 8346: data <= 'd0; 8347: data <= 'd0; 8348: data <= 'd0; 8349: data <= 'd0; 8350: data <= 'd0; 8351: data <= 'd0; 8352: data <= 'd0; 8353: data <= 'd0; 8354: data <= 'd0; 8355: data <= 'd0; 8356: data <= 'd0; 8357: data <= 'd0; 8358: data <= 'd0; 8359: data <= 'd0; 8360: data <= 'd0; 8361: data <= 'd0; 8362: data <= 'd0; 8363: data <= 'd0; 8364: data <= 'd0; 8365: data <= 'd0; 8366: data <= 'd0; 8367: data <= 'd0; 8368: data <= 'd0; 8369: data <= 'd0; 8370: data <= 'd0; 8371: data <= 'd0; 8372: data <= 'd0; 8373: data <= 'd0; 8374: data <= 'd0; 8375: data <= 'd0; 8376: data <= 'd0; 8377: data <= 'd0; 8378: data <= 'd0; 8379: data <= 'd0; 8380: data <= 'd0; 8381: data <= 'd0; 8382: data <= 'd0; 8383: data <= 'd0; 8384: data <= 'd0; 8385: data <= 'd0; 8386: data <= 'd0; 8387: data <= 'd0; 8388: data <= 'd0; 8389: data <= 'd0; 8390: data <= 'd0; 8391: data <= 'd0; 8392: data <= 'd0; 8393: data <= 'd0; 8394: data <= 'd0; 8395: data <= 'd0; 8396: data <= 'd0; 8397: data <= 'd0; 8398: data <= 'd0; 8399: data <= 'd0; 8400: data <= 'd0; 8401: data <= 'd0; 8402: data <= 'd0; 8403: data <= 'd0; 8404: data <= 'd0; 8405: data <= 'd0; 8406: data <= 'd0; 8407: data <= 'd0; 8408: data <= 'd0; 8409: data <= 'd0; 8410: data <= 'd0; 8411: data <= 'd0; 8412: data <= 'd0; 8413: data <= 'd0; 8414: data <= 'd0; 8415: data <= 'd0; 8416: data <= 'd0; 8417: data <= 'd0; 8418: data <= 'd0; 8419: data <= 'd0; 8420: data <= 'd0; 8421: data <= 'd0; 8422: data <= 'd0; 8423: data <= 'd0; 8424: data <= 'd0; 8425: data <= 'd0; 8426: data <= 'd0; 8427: data <= 'd0; 8428: data <= 'd0; 8429: data <= 'd0; 8430: data <= 'd0; 8431: data <= 'd0; 8432: data <= 'd0; 8433: data <= 'd0; 8434: data <= 'd0; 8435: data <= 'd0; 8436: data <= 'd0; 8437: data <= 'd0; 8438: data <= 'd0; 8439: data <= 'd0; 8440: data <= 'd0; 8441: data <= 'd0; 8442: data <= 'd0; 8443: data <= 'd0; 8444: data <= 'd0; 8445: data <= 'd0; 8446: data <= 'd0; 8447: data <= 'd0; 8448: data <= 'd0; 8449: data <= 'd0; 8450: data <= 'd0; 8451: data <= 'd0; 8452: data <= 'd0; 8453: data <= 'd0; 8454: data <= 'd0; 8455: data <= 'd0; 8456: data <= 'd0; 8457: data <= 'd0; 8458: data <= 'd0; 8459: data <= 'd0; 8460: data <= 'd0; 8461: data <= 'd0; 8462: data <= 'd0; 8463: data <= 'd0; 8464: data <= 'd0; 8465: data <= 'd0; 8466: data <= 'd0; 8467: data <= 'd0; 8468: data <= 'd0; 8469: data <= 'd0; 8470: data <= 'd0; 8471: data <= 'd0; 8472: data <= 'd0; 8473: data <= 'd0; 8474: data <= 'd0; 8475: data <= 'd0; 8476: data <= 'd0; 8477: data <= 'd0; 8478: data <= 'd0; 8479: data <= 'd0; 8480: data <= 'd0; 8481: data <= 'd0; 8482: data <= 'd0; 8483: data <= 'd0; 8484: data <= 'd0; 8485: data <= 'd0; 8486: data <= 'd0; 8487: data <= 'd0; 8488: data <= 'd0; 8489: data <= 'd0; 8490: data <= 'd0; 8491: data <= 'd0; 8492: data <= 'd2; 8493: data <= 'd2; 8494: data <= 'd2; 8495: data <= 'd2; 8496: data <= 'd2; 8497: data <= 'd2; 8498: data <= 'd0; 8499: data <= 'd0; 8500: data <= 'd0; 8501: data <= 'd0; 8502: data <= 'd0; 8503: data <= 'd0; 8504: data <= 'd0; 8505: data <= 'd0; 8506: data <= 'd0; 8507: data <= 'd0; 8508: data <= 'd0; 8509: data <= 'd0; 8510: data <= 'd0; 8511: data <= 'd0; 8512: data <= 'd0; 8513: data <= 'd0; 8514: data <= 'd0; 8515: data <= 'd0; 8516: data <= 'd0; 8517: data <= 'd0; 8518: data <= 'd0; 8519: data <= 'd0; 8520: data <= 'd0; 8521: data <= 'd0; 8522: data <= 'd2; 8523: data <= 'd2; 8524: data <= 'd6; 8525: data <= 'd6; 8526: data <= 'd6; 8527: data <= 'd6; 8528: data <= 'd6; 8529: data <= 'd6; 8530: data <= 'd2; 8531: data <= 'd2; 8532: data <= 'd0; 8533: data <= 'd0; 8534: data <= 'd0; 8535: data <= 'd0; 8536: data <= 'd0; 8537: data <= 'd0; 8538: data <= 'd0; 8539: data <= 'd0; 8540: data <= 'd0; 8541: data <= 'd0; 8542: data <= 'd0; 8543: data <= 'd0; 8544: data <= 'd0; 8545: data <= 'd0; 8546: data <= 'd0; 8547: data <= 'd0; 8548: data <= 'd0; 8549: data <= 'd0; 8550: data <= 'd0; 8551: data <= 'd0; 8552: data <= 'd0; 8553: data <= 'd2; 8554: data <= 'd1; 8555: data <= 'd3; 8556: data <= 'd6; 8557: data <= 'd6; 8558: data <= 'd6; 8559: data <= 'd6; 8560: data <= 'd6; 8561: data <= 'd6; 8562: data <= 'd6; 8563: data <= 'd3; 8564: data <= 'd2; 8565: data <= 'd0; 8566: data <= 'd0; 8567: data <= 'd0; 8568: data <= 'd0; 8569: data <= 'd0; 8570: data <= 'd0; 8571: data <= 'd0; 8572: data <= 'd0; 8573: data <= 'd0; 8574: data <= 'd0; 8575: data <= 'd0; 8576: data <= 'd0; 8577: data <= 'd0; 8578: data <= 'd0; 8579: data <= 'd0; 8580: data <= 'd0; 8581: data <= 'd0; 8582: data <= 'd0; 8583: data <= 'd0; 8584: data <= 'd2; 8585: data <= 'd1; 8586: data <= 'd1; 8587: data <= 'd1; 8588: data <= 'd3; 8589: data <= 'd6; 8590: data <= 'd6; 8591: data <= 'd6; 8592: data <= 'd6; 8593: data <= 'd6; 8594: data <= 'd3; 8595: data <= 'd1; 8596: data <= 'd1; 8597: data <= 'd2; 8598: data <= 'd0; 8599: data <= 'd0; 8600: data <= 'd0; 8601: data <= 'd0; 8602: data <= 'd0; 8603: data <= 'd0; 8604: data <= 'd0; 8605: data <= 'd0; 8606: data <= 'd0; 8607: data <= 'd0; 8608: data <= 'd0; 8609: data <= 'd0; 8610: data <= 'd0; 8611: data <= 'd0; 8612: data <= 'd0; 8613: data <= 'd0; 8614: data <= 'd0; 8615: data <= 'd0; 8616: data <= 'd2; 8617: data <= 'd1; 8618: data <= 'd1; 8619: data <= 'd5; 8620: data <= 'd5; 8621: data <= 'd5; 8622: data <= 'd1; 8623: data <= 'd1; 8624: data <= 'd1; 8625: data <= 'd1; 8626: data <= 'd1; 8627: data <= 'd5; 8628: data <= 'd5; 8629: data <= 'd2; 8630: data <= 'd0; 8631: data <= 'd0; 8632: data <= 'd0; 8633: data <= 'd0; 8634: data <= 'd0; 8635: data <= 'd0; 8636: data <= 'd0; 8637: data <= 'd0; 8638: data <= 'd0; 8639: data <= 'd0; 8640: data <= 'd0; 8641: data <= 'd0; 8642: data <= 'd0; 8643: data <= 'd0; 8644: data <= 'd0; 8645: data <= 'd0; 8646: data <= 'd0; 8647: data <= 'd2; 8648: data <= 'd1; 8649: data <= 'd5; 8650: data <= 'd5; 8651: data <= 'd3; 8652: data <= 'd6; 8653: data <= 'd6; 8654: data <= 'd6; 8655: data <= 'd6; 8656: data <= 'd6; 8657: data <= 'd6; 8658: data <= 'd6; 8659: data <= 'd6; 8660: data <= 'd3; 8661: data <= 'd5; 8662: data <= 'd2; 8663: data <= 'd0; 8664: data <= 'd0; 8665: data <= 'd0; 8666: data <= 'd0; 8667: data <= 'd0; 8668: data <= 'd0; 8669: data <= 'd0; 8670: data <= 'd0; 8671: data <= 'd0; 8672: data <= 'd0; 8673: data <= 'd0; 8674: data <= 'd0; 8675: data <= 'd0; 8676: data <= 'd0; 8677: data <= 'd0; 8678: data <= 'd0; 8679: data <= 'd2; 8680: data <= 'd5; 8681: data <= 'd3; 8682: data <= 'd6; 8683: data <= 'd3; 8684: data <= 'd1; 8685: data <= 'd1; 8686: data <= 'd1; 8687: data <= 'd1; 8688: data <= 'd1; 8689: data <= 'd1; 8690: data <= 'd1; 8691: data <= 'd1; 8692: data <= 'd1; 8693: data <= 'd3; 8694: data <= 'd2; 8695: data <= 'd0; 8696: data <= 'd0; 8697: data <= 'd0; 8698: data <= 'd0; 8699: data <= 'd0; 8700: data <= 'd0; 8701: data <= 'd0; 8702: data <= 'd0; 8703: data <= 'd0; 8704: data <= 'd0; 8705: data <= 'd0; 8706: data <= 'd0; 8707: data <= 'd0; 8708: data <= 'd0; 8709: data <= 'd0; 8710: data <= 'd0; 8711: data <= 'd2; 8712: data <= 'd5; 8713: data <= 'd3; 8714: data <= 'd1; 8715: data <= 'd1; 8716: data <= 'd1; 8717: data <= 'd5; 8718: data <= 'd5; 8719: data <= 'd5; 8720: data <= 'd5; 8721: data <= 'd5; 8722: data <= 'd5; 8723: data <= 'd5; 8724: data <= 'd1; 8725: data <= 'd1; 8726: data <= 'd2; 8727: data <= 'd0; 8728: data <= 'd0; 8729: data <= 'd0; 8730: data <= 'd0; 8731: data <= 'd0; 8732: data <= 'd0; 8733: data <= 'd0; 8734: data <= 'd0; 8735: data <= 'd0; 8736: data <= 'd0; 8737: data <= 'd0; 8738: data <= 'd0; 8739: data <= 'd0; 8740: data <= 'd0; 8741: data <= 'd0; 8742: data <= 'd0; 8743: data <= 'd2; 8744: data <= 'd6; 8745: data <= 'd1; 8746: data <= 'd5; 8747: data <= 'd2; 8748: data <= 'd2; 8749: data <= 'd2; 8750: data <= 'd2; 8751: data <= 'd2; 8752: data <= 'd2; 8753: data <= 'd2; 8754: data <= 'd2; 8755: data <= 'd2; 8756: data <= 'd2; 8757: data <= 'd5; 8758: data <= 'd2; 8759: data <= 'd0; 8760: data <= 'd0; 8761: data <= 'd0; 8762: data <= 'd0; 8763: data <= 'd0; 8764: data <= 'd0; 8765: data <= 'd0; 8766: data <= 'd0; 8767: data <= 'd0; 8768: data <= 'd0; 8769: data <= 'd0; 8770: data <= 'd0; 8771: data <= 'd0; 8772: data <= 'd0; 8773: data <= 'd2; 8774: data <= 'd2; 8775: data <= 'd2; 8776: data <= 'd1; 8777: data <= 'd5; 8778: data <= 'd2; 8779: data <= 'd8; 8780: data <= 'd8; 8781: data <= 'd8; 8782: data <= 'd8; 8783: data <= 'd8; 8784: data <= 'd9; 8785: data <= 'd9; 8786: data <= 'd8; 8787: data <= 'd8; 8788: data <= 'd8; 8789: data <= 'd2; 8790: data <= 'd2; 8791: data <= 'd0; 8792: data <= 'd0; 8793: data <= 'd0; 8794: data <= 'd0; 8795: data <= 'd0; 8796: data <= 'd0; 8797: data <= 'd0; 8798: data <= 'd0; 8799: data <= 'd0; 8800: data <= 'd0; 8801: data <= 'd0; 8802: data <= 'd0; 8803: data <= 'd0; 8804: data <= 'd0; 8805: data <= 'd2; 8806: data <= 'd1; 8807: data <= 'd2; 8808: data <= 'd1; 8809: data <= 'd2; 8810: data <= 'd8; 8811: data <= 'd8; 8812: data <= 'd9; 8813: data <= 'd9; 8814: data <= 'd2; 8815: data <= 'd9; 8816: data <= 'd11; 8817: data <= 'd11; 8818: data <= 'd10; 8819: data <= 'd2; 8820: data <= 'd9; 8821: data <= 'd2; 8822: data <= 'd2; 8823: data <= 'd0; 8824: data <= 'd0; 8825: data <= 'd0; 8826: data <= 'd0; 8827: data <= 'd0; 8828: data <= 'd0; 8829: data <= 'd0; 8830: data <= 'd0; 8831: data <= 'd0; 8832: data <= 'd0; 8833: data <= 'd0; 8834: data <= 'd0; 8835: data <= 'd0; 8836: data <= 'd0; 8837: data <= 'd2; 8838: data <= 'd5; 8839: data <= 'd1; 8840: data <= 'd2; 8841: data <= 'd9; 8842: data <= 'd10; 8843: data <= 'd9; 8844: data <= 'd9; 8845: data <= 'd10; 8846: data <= 'd11; 8847: data <= 'd10; 8848: data <= 'd11; 8849: data <= 'd11; 8850: data <= 'd10; 8851: data <= 'd11; 8852: data <= 'd10; 8853: data <= 'd9; 8854: data <= 'd2; 8855: data <= 'd0; 8856: data <= 'd0; 8857: data <= 'd0; 8858: data <= 'd0; 8859: data <= 'd0; 8860: data <= 'd0; 8861: data <= 'd0; 8862: data <= 'd0; 8863: data <= 'd0; 8864: data <= 'd0; 8865: data <= 'd0; 8866: data <= 'd0; 8867: data <= 'd0; 8868: data <= 'd0; 8869: data <= 'd0; 8870: data <= 'd2; 8871: data <= 'd5; 8872: data <= 'd5; 8873: data <= 'd2; 8874: data <= 'd8; 8875: data <= 'd9; 8876: data <= 'd9; 8877: data <= 'd10; 8878: data <= 'd10; 8879: data <= 'd10; 8880: data <= 'd8; 8881: data <= 'd8; 8882: data <= 'd10; 8883: data <= 'd10; 8884: data <= 'd9; 8885: data <= 'd2; 8886: data <= 'd0; 8887: data <= 'd0; 8888: data <= 'd0; 8889: data <= 'd0; 8890: data <= 'd0; 8891: data <= 'd0; 8892: data <= 'd0; 8893: data <= 'd0; 8894: data <= 'd0; 8895: data <= 'd0; 8896: data <= 'd0; 8897: data <= 'd0; 8898: data <= 'd0; 8899: data <= 'd0; 8900: data <= 'd0; 8901: data <= 'd0; 8902: data <= 'd0; 8903: data <= 'd2; 8904: data <= 'd2; 8905: data <= 'd2; 8906: data <= 'd8; 8907: data <= 'd8; 8908: data <= 'd9; 8909: data <= 'd9; 8910: data <= 'd10; 8911: data <= 'd10; 8912: data <= 'd9; 8913: data <= 'd9; 8914: data <= 'd10; 8915: data <= 'd10; 8916: data <= 'd9; 8917: data <= 'd2; 8918: data <= 'd0; 8919: data <= 'd0; 8920: data <= 'd0; 8921: data <= 'd0; 8922: data <= 'd0; 8923: data <= 'd0; 8924: data <= 'd0; 8925: data <= 'd0; 8926: data <= 'd0; 8927: data <= 'd0; 8928: data <= 'd0; 8929: data <= 'd0; 8930: data <= 'd0; 8931: data <= 'd0; 8932: data <= 'd0; 8933: data <= 'd0; 8934: data <= 'd0; 8935: data <= 'd0; 8936: data <= 'd0; 8937: data <= 'd2; 8938: data <= 'd2; 8939: data <= 'd5; 8940: data <= 'd5; 8941: data <= 'd8; 8942: data <= 'd9; 8943: data <= 'd9; 8944: data <= 'd9; 8945: data <= 'd9; 8946: data <= 'd9; 8947: data <= 'd9; 8948: data <= 'd5; 8949: data <= 'd2; 8950: data <= 'd0; 8951: data <= 'd0; 8952: data <= 'd0; 8953: data <= 'd0; 8954: data <= 'd0; 8955: data <= 'd0; 8956: data <= 'd0; 8957: data <= 'd0; 8958: data <= 'd0; 8959: data <= 'd0; 8960: data <= 'd0; 8961: data <= 'd0; 8962: data <= 'd0; 8963: data <= 'd0; 8964: data <= 'd0; 8965: data <= 'd0; 8966: data <= 'd0; 8967: data <= 'd0; 8968: data <= 'd2; 8969: data <= 'd7; 8970: data <= 'd1; 8971: data <= 'd1; 8972: data <= 'd1; 8973: data <= 'd3; 8974: data <= 'd3; 8975: data <= 'd3; 8976: data <= 'd5; 8977: data <= 'd5; 8978: data <= 'd3; 8979: data <= 'd3; 8980: data <= 'd1; 8981: data <= 'd2; 8982: data <= 'd0; 8983: data <= 'd0; 8984: data <= 'd0; 8985: data <= 'd0; 8986: data <= 'd0; 8987: data <= 'd0; 8988: data <= 'd0; 8989: data <= 'd0; 8990: data <= 'd0; 8991: data <= 'd0; 8992: data <= 'd0; 8993: data <= 'd0; 8994: data <= 'd0; 8995: data <= 'd0; 8996: data <= 'd0; 8997: data <= 'd0; 8998: data <= 'd0; 8999: data <= 'd0; 9000: data <= 'd2; 9001: data <= 'd7; 9002: data <= 'd7; 9003: data <= 'd5; 9004: data <= 'd1; 9005: data <= 'd3; 9006: data <= 'd3; 9007: data <= 'd3; 9008: data <= 'd1; 9009: data <= 'd1; 9010: data <= 'd3; 9011: data <= 'd3; 9012: data <= 'd1; 9013: data <= 'd2; 9014: data <= 'd2; 9015: data <= 'd0; 9016: data <= 'd0; 9017: data <= 'd0; 9018: data <= 'd0; 9019: data <= 'd0; 9020: data <= 'd0; 9021: data <= 'd0; 9022: data <= 'd0; 9023: data <= 'd0; 9024: data <= 'd0; 9025: data <= 'd0; 9026: data <= 'd0; 9027: data <= 'd0; 9028: data <= 'd0; 9029: data <= 'd0; 9030: data <= 'd0; 9031: data <= 'd0; 9032: data <= 'd0; 9033: data <= 'd2; 9034: data <= 'd9; 9035: data <= 'd9; 9036: data <= 'd2; 9037: data <= 'd1; 9038: data <= 'd3; 9039: data <= 'd3; 9040: data <= 'd1; 9041: data <= 'd1; 9042: data <= 'd3; 9043: data <= 'd1; 9044: data <= 'd1; 9045: data <= 'd8; 9046: data <= 'd9; 9047: data <= 'd2; 9048: data <= 'd0; 9049: data <= 'd0; 9050: data <= 'd0; 9051: data <= 'd0; 9052: data <= 'd0; 9053: data <= 'd0; 9054: data <= 'd0; 9055: data <= 'd0; 9056: data <= 'd0; 9057: data <= 'd0; 9058: data <= 'd0; 9059: data <= 'd0; 9060: data <= 'd0; 9061: data <= 'd0; 9062: data <= 'd0; 9063: data <= 'd0; 9064: data <= 'd0; 9065: data <= 'd2; 9066: data <= 'd9; 9067: data <= 'd9; 9068: data <= 'd2; 9069: data <= 'd2; 9070: data <= 'd2; 9071: data <= 'd5; 9072: data <= 'd5; 9073: data <= 'd5; 9074: data <= 'd2; 9075: data <= 'd2; 9076: data <= 'd2; 9077: data <= 'd8; 9078: data <= 'd9; 9079: data <= 'd2; 9080: data <= 'd0; 9081: data <= 'd0; 9082: data <= 'd0; 9083: data <= 'd0; 9084: data <= 'd0; 9085: data <= 'd0; 9086: data <= 'd0; 9087: data <= 'd0; 9088: data <= 'd0; 9089: data <= 'd0; 9090: data <= 'd0; 9091: data <= 'd0; 9092: data <= 'd0; 9093: data <= 'd0; 9094: data <= 'd0; 9095: data <= 'd0; 9096: data <= 'd0; 9097: data <= 'd0; 9098: data <= 'd2; 9099: data <= 'd2; 9100: data <= 'd1; 9101: data <= 'd3; 9102: data <= 'd3; 9103: data <= 'd3; 9104: data <= 'd1; 9105: data <= 'd3; 9106: data <= 'd3; 9107: data <= 'd3; 9108: data <= 'd2; 9109: data <= 'd2; 9110: data <= 'd2; 9111: data <= 'd0; 9112: data <= 'd0; 9113: data <= 'd0; 9114: data <= 'd0; 9115: data <= 'd0; 9116: data <= 'd0; 9117: data <= 'd0; 9118: data <= 'd0; 9119: data <= 'd0; 9120: data <= 'd0; 9121: data <= 'd0; 9122: data <= 'd0; 9123: data <= 'd0; 9124: data <= 'd0; 9125: data <= 'd0; 9126: data <= 'd0; 9127: data <= 'd0; 9128: data <= 'd0; 9129: data <= 'd0; 9130: data <= 'd2; 9131: data <= 'd4; 9132: data <= 'd7; 9133: data <= 'd7; 9134: data <= 'd2; 9135: data <= 'd2; 9136: data <= 'd2; 9137: data <= 'd5; 9138: data <= 'd5; 9139: data <= 'd4; 9140: data <= 'd2; 9141: data <= 'd0; 9142: data <= 'd0; 9143: data <= 'd0; 9144: data <= 'd0; 9145: data <= 'd0; 9146: data <= 'd0; 9147: data <= 'd0; 9148: data <= 'd0; 9149: data <= 'd0; 9150: data <= 'd0; 9151: data <= 'd0; 9152: data <= 'd0; 9153: data <= 'd0; 9154: data <= 'd0; 9155: data <= 'd0; 9156: data <= 'd0; 9157: data <= 'd0; 9158: data <= 'd0; 9159: data <= 'd0; 9160: data <= 'd0; 9161: data <= 'd0; 9162: data <= 'd0; 9163: data <= 'd2; 9164: data <= 'd4; 9165: data <= 'd7; 9166: data <= 'd2; 9167: data <= 'd0; 9168: data <= 'd0; 9169: data <= 'd2; 9170: data <= 'd4; 9171: data <= 'd4; 9172: data <= 'd2; 9173: data <= 'd0; 9174: data <= 'd0; 9175: data <= 'd0; 9176: data <= 'd0; 9177: data <= 'd0; 9178: data <= 'd0; 9179: data <= 'd0; 9180: data <= 'd0; 9181: data <= 'd0; 9182: data <= 'd0; 9183: data <= 'd0; 9184: data <= 'd0; 9185: data <= 'd0; 9186: data <= 'd0; 9187: data <= 'd0; 9188: data <= 'd0; 9189: data <= 'd0; 9190: data <= 'd0; 9191: data <= 'd0; 9192: data <= 'd0; 9193: data <= 'd0; 9194: data <= 'd0; 9195: data <= 'd2; 9196: data <= 'd2; 9197: data <= 'd2; 9198: data <= 'd2; 9199: data <= 'd0; 9200: data <= 'd0; 9201: data <= 'd0; 9202: data <= 'd2; 9203: data <= 'd2; 9204: data <= 'd2; 9205: data <= 'd0; 9206: data <= 'd0; 9207: data <= 'd0; 9208: data <= 'd0; 9209: data <= 'd0; 9210: data <= 'd0; 9211: data <= 'd0; 9212: data <= 'd0; 9213: data <= 'd0; 9214: data <= 'd0; 9215: data <= 'd0; 9216: data <= 'd0; 9217: data <= 'd0; 9218: data <= 'd0; 9219: data <= 'd0; 9220: data <= 'd0; 9221: data <= 'd0; 9222: data <= 'd0; 9223: data <= 'd0; 9224: data <= 'd0; 9225: data <= 'd0; 9226: data <= 'd0; 9227: data <= 'd0; 9228: data <= 'd0; 9229: data <= 'd0; 9230: data <= 'd0; 9231: data <= 'd0; 9232: data <= 'd0; 9233: data <= 'd0; 9234: data <= 'd0; 9235: data <= 'd0; 9236: data <= 'd0; 9237: data <= 'd0; 9238: data <= 'd0; 9239: data <= 'd0; 9240: data <= 'd0; 9241: data <= 'd0; 9242: data <= 'd0; 9243: data <= 'd0; 9244: data <= 'd0; 9245: data <= 'd0; 9246: data <= 'd0; 9247: data <= 'd0; 9248: data <= 'd0; 9249: data <= 'd0; 9250: data <= 'd0; 9251: data <= 'd0; 9252: data <= 'd0; 9253: data <= 'd0; 9254: data <= 'd0; 9255: data <= 'd0; 9256: data <= 'd0; 9257: data <= 'd0; 9258: data <= 'd0; 9259: data <= 'd0; 9260: data <= 'd0; 9261: data <= 'd0; 9262: data <= 'd0; 9263: data <= 'd0; 9264: data <= 'd0; 9265: data <= 'd0; 9266: data <= 'd0; 9267: data <= 'd0; 9268: data <= 'd0; 9269: data <= 'd0; 9270: data <= 'd0; 9271: data <= 'd0; 9272: data <= 'd0; 9273: data <= 'd0; 9274: data <= 'd0; 9275: data <= 'd0; 9276: data <= 'd0; 9277: data <= 'd0; 9278: data <= 'd0; 9279: data <= 'd0; 9280: data <= 'd0; 9281: data <= 'd0; 9282: data <= 'd0; 9283: data <= 'd0; 9284: data <= 'd0; 9285: data <= 'd0; 9286: data <= 'd0; 9287: data <= 'd0; 9288: data <= 'd0; 9289: data <= 'd0; 9290: data <= 'd0; 9291: data <= 'd0; 9292: data <= 'd0; 9293: data <= 'd0; 9294: data <= 'd0; 9295: data <= 'd0; 9296: data <= 'd0; 9297: data <= 'd0; 9298: data <= 'd0; 9299: data <= 'd0; 9300: data <= 'd0; 9301: data <= 'd0; 9302: data <= 'd0; 9303: data <= 'd0; 9304: data <= 'd0; 9305: data <= 'd0; 9306: data <= 'd0; 9307: data <= 'd0; 9308: data <= 'd0; 9309: data <= 'd0; 9310: data <= 'd0; 9311: data <= 'd0; 9312: data <= 'd0; 9313: data <= 'd0; 9314: data <= 'd0; 9315: data <= 'd0; 9316: data <= 'd0; 9317: data <= 'd0; 9318: data <= 'd0; 9319: data <= 'd0; 9320: data <= 'd0; 9321: data <= 'd0; 9322: data <= 'd0; 9323: data <= 'd0; 9324: data <= 'd0; 9325: data <= 'd0; 9326: data <= 'd0; 9327: data <= 'd0; 9328: data <= 'd0; 9329: data <= 'd0; 9330: data <= 'd0; 9331: data <= 'd0; 9332: data <= 'd0; 9333: data <= 'd0; 9334: data <= 'd0; 9335: data <= 'd0; 9336: data <= 'd0; 9337: data <= 'd0; 9338: data <= 'd0; 9339: data <= 'd0; 9340: data <= 'd0; 9341: data <= 'd0; 9342: data <= 'd0; 9343: data <= 'd0; 9344: data <= 'd0; 9345: data <= 'd0; 9346: data <= 'd0; 9347: data <= 'd0; 9348: data <= 'd0; 9349: data <= 'd0; 9350: data <= 'd0; 9351: data <= 'd0; 9352: data <= 'd0; 9353: data <= 'd0; 9354: data <= 'd0; 9355: data <= 'd0; 9356: data <= 'd0; 9357: data <= 'd0; 9358: data <= 'd0; 9359: data <= 'd0; 9360: data <= 'd0; 9361: data <= 'd0; 9362: data <= 'd0; 9363: data <= 'd0; 9364: data <= 'd0; 9365: data <= 'd0; 9366: data <= 'd0; 9367: data <= 'd0; 9368: data <= 'd0; 9369: data <= 'd0; 9370: data <= 'd0; 9371: data <= 'd0; 9372: data <= 'd0; 9373: data <= 'd0; 9374: data <= 'd0; 9375: data <= 'd0; 9376: data <= 'd0; 9377: data <= 'd0; 9378: data <= 'd0; 9379: data <= 'd0; 9380: data <= 'd0; 9381: data <= 'd0; 9382: data <= 'd0; 9383: data <= 'd0; 9384: data <= 'd0; 9385: data <= 'd0; 9386: data <= 'd0; 9387: data <= 'd0; 9388: data <= 'd0; 9389: data <= 'd0; 9390: data <= 'd0; 9391: data <= 'd0; 9392: data <= 'd0; 9393: data <= 'd0; 9394: data <= 'd0; 9395: data <= 'd0; 9396: data <= 'd0; 9397: data <= 'd0; 9398: data <= 'd0; 9399: data <= 'd0; 9400: data <= 'd0; 9401: data <= 'd0; 9402: data <= 'd0; 9403: data <= 'd0; 9404: data <= 'd0; 9405: data <= 'd0; 9406: data <= 'd0; 9407: data <= 'd0; 9408: data <= 'd0; 9409: data <= 'd0; 9410: data <= 'd0; 9411: data <= 'd0; 9412: data <= 'd0; 9413: data <= 'd0; 9414: data <= 'd0; 9415: data <= 'd0; 9416: data <= 'd0; 9417: data <= 'd0; 9418: data <= 'd0; 9419: data <= 'd0; 9420: data <= 'd0; 9421: data <= 'd0; 9422: data <= 'd0; 9423: data <= 'd0; 9424: data <= 'd0; 9425: data <= 'd0; 9426: data <= 'd0; 9427: data <= 'd0; 9428: data <= 'd0; 9429: data <= 'd0; 9430: data <= 'd0; 9431: data <= 'd0; 9432: data <= 'd0; 9433: data <= 'd0; 9434: data <= 'd0; 9435: data <= 'd0; 9436: data <= 'd0; 9437: data <= 'd0; 9438: data <= 'd0; 9439: data <= 'd0; 9440: data <= 'd0; 9441: data <= 'd0; 9442: data <= 'd0; 9443: data <= 'd0; 9444: data <= 'd0; 9445: data <= 'd0; 9446: data <= 'd0; 9447: data <= 'd0; 9448: data <= 'd0; 9449: data <= 'd0; 9450: data <= 'd0; 9451: data <= 'd0; 9452: data <= 'd0; 9453: data <= 'd0; 9454: data <= 'd0; 9455: data <= 'd0; 9456: data <= 'd0; 9457: data <= 'd0; 9458: data <= 'd0; 9459: data <= 'd0; 9460: data <= 'd0; 9461: data <= 'd0; 9462: data <= 'd0; 9463: data <= 'd0; 9464: data <= 'd0; 9465: data <= 'd0; 9466: data <= 'd0; 9467: data <= 'd0; 9468: data <= 'd0; 9469: data <= 'd0; 9470: data <= 'd0; 9471: data <= 'd0; 9472: data <= 'd0; 9473: data <= 'd0; 9474: data <= 'd0; 9475: data <= 'd0; 9476: data <= 'd0; 9477: data <= 'd0; 9478: data <= 'd0; 9479: data <= 'd0; 9480: data <= 'd0; 9481: data <= 'd0; 9482: data <= 'd0; 9483: data <= 'd0; 9484: data <= 'd0; 9485: data <= 'd0; 9486: data <= 'd0; 9487: data <= 'd0; 9488: data <= 'd0; 9489: data <= 'd0; 9490: data <= 'd0; 9491: data <= 'd0; 9492: data <= 'd0; 9493: data <= 'd0; 9494: data <= 'd0; 9495: data <= 'd0; 9496: data <= 'd0; 9497: data <= 'd0; 9498: data <= 'd0; 9499: data <= 'd0; 9500: data <= 'd0; 9501: data <= 'd0; 9502: data <= 'd0; 9503: data <= 'd0; 9504: data <= 'd0; 9505: data <= 'd0; 9506: data <= 'd0; 9507: data <= 'd0; 9508: data <= 'd0; 9509: data <= 'd0; 9510: data <= 'd0; 9511: data <= 'd0; 9512: data <= 'd0; 9513: data <= 'd0; 9514: data <= 'd2; 9515: data <= 'd2; 9516: data <= 'd2; 9517: data <= 'd2; 9518: data <= 'd2; 9519: data <= 'd2; 9520: data <= 'd0; 9521: data <= 'd0; 9522: data <= 'd0; 9523: data <= 'd0; 9524: data <= 'd0; 9525: data <= 'd0; 9526: data <= 'd0; 9527: data <= 'd0; 9528: data <= 'd0; 9529: data <= 'd0; 9530: data <= 'd0; 9531: data <= 'd0; 9532: data <= 'd0; 9533: data <= 'd0; 9534: data <= 'd0; 9535: data <= 'd0; 9536: data <= 'd0; 9537: data <= 'd0; 9538: data <= 'd0; 9539: data <= 'd0; 9540: data <= 'd0; 9541: data <= 'd0; 9542: data <= 'd0; 9543: data <= 'd0; 9544: data <= 'd2; 9545: data <= 'd2; 9546: data <= 'd6; 9547: data <= 'd6; 9548: data <= 'd6; 9549: data <= 'd6; 9550: data <= 'd6; 9551: data <= 'd6; 9552: data <= 'd2; 9553: data <= 'd2; 9554: data <= 'd0; 9555: data <= 'd0; 9556: data <= 'd0; 9557: data <= 'd0; 9558: data <= 'd0; 9559: data <= 'd0; 9560: data <= 'd0; 9561: data <= 'd0; 9562: data <= 'd0; 9563: data <= 'd0; 9564: data <= 'd0; 9565: data <= 'd0; 9566: data <= 'd0; 9567: data <= 'd0; 9568: data <= 'd0; 9569: data <= 'd0; 9570: data <= 'd0; 9571: data <= 'd0; 9572: data <= 'd0; 9573: data <= 'd0; 9574: data <= 'd0; 9575: data <= 'd2; 9576: data <= 'd1; 9577: data <= 'd3; 9578: data <= 'd6; 9579: data <= 'd6; 9580: data <= 'd6; 9581: data <= 'd6; 9582: data <= 'd6; 9583: data <= 'd6; 9584: data <= 'd6; 9585: data <= 'd3; 9586: data <= 'd2; 9587: data <= 'd0; 9588: data <= 'd0; 9589: data <= 'd0; 9590: data <= 'd0; 9591: data <= 'd0; 9592: data <= 'd0; 9593: data <= 'd0; 9594: data <= 'd0; 9595: data <= 'd0; 9596: data <= 'd0; 9597: data <= 'd0; 9598: data <= 'd0; 9599: data <= 'd0; 9600: data <= 'd0; 9601: data <= 'd0; 9602: data <= 'd0; 9603: data <= 'd0; 9604: data <= 'd0; 9605: data <= 'd0; 9606: data <= 'd2; 9607: data <= 'd1; 9608: data <= 'd1; 9609: data <= 'd1; 9610: data <= 'd3; 9611: data <= 'd6; 9612: data <= 'd6; 9613: data <= 'd6; 9614: data <= 'd6; 9615: data <= 'd6; 9616: data <= 'd3; 9617: data <= 'd1; 9618: data <= 'd1; 9619: data <= 'd2; 9620: data <= 'd0; 9621: data <= 'd0; 9622: data <= 'd0; 9623: data <= 'd0; 9624: data <= 'd0; 9625: data <= 'd0; 9626: data <= 'd0; 9627: data <= 'd0; 9628: data <= 'd0; 9629: data <= 'd0; 9630: data <= 'd0; 9631: data <= 'd0; 9632: data <= 'd0; 9633: data <= 'd0; 9634: data <= 'd0; 9635: data <= 'd0; 9636: data <= 'd0; 9637: data <= 'd0; 9638: data <= 'd2; 9639: data <= 'd1; 9640: data <= 'd1; 9641: data <= 'd5; 9642: data <= 'd5; 9643: data <= 'd5; 9644: data <= 'd1; 9645: data <= 'd1; 9646: data <= 'd1; 9647: data <= 'd1; 9648: data <= 'd1; 9649: data <= 'd5; 9650: data <= 'd5; 9651: data <= 'd2; 9652: data <= 'd0; 9653: data <= 'd0; 9654: data <= 'd0; 9655: data <= 'd0; 9656: data <= 'd0; 9657: data <= 'd0; 9658: data <= 'd0; 9659: data <= 'd0; 9660: data <= 'd0; 9661: data <= 'd0; 9662: data <= 'd0; 9663: data <= 'd0; 9664: data <= 'd0; 9665: data <= 'd0; 9666: data <= 'd0; 9667: data <= 'd0; 9668: data <= 'd0; 9669: data <= 'd2; 9670: data <= 'd1; 9671: data <= 'd5; 9672: data <= 'd5; 9673: data <= 'd3; 9674: data <= 'd6; 9675: data <= 'd6; 9676: data <= 'd6; 9677: data <= 'd6; 9678: data <= 'd6; 9679: data <= 'd6; 9680: data <= 'd6; 9681: data <= 'd6; 9682: data <= 'd3; 9683: data <= 'd5; 9684: data <= 'd2; 9685: data <= 'd0; 9686: data <= 'd0; 9687: data <= 'd0; 9688: data <= 'd0; 9689: data <= 'd0; 9690: data <= 'd0; 9691: data <= 'd0; 9692: data <= 'd0; 9693: data <= 'd0; 9694: data <= 'd0; 9695: data <= 'd0; 9696: data <= 'd0; 9697: data <= 'd0; 9698: data <= 'd0; 9699: data <= 'd0; 9700: data <= 'd0; 9701: data <= 'd2; 9702: data <= 'd5; 9703: data <= 'd3; 9704: data <= 'd6; 9705: data <= 'd3; 9706: data <= 'd1; 9707: data <= 'd1; 9708: data <= 'd1; 9709: data <= 'd1; 9710: data <= 'd1; 9711: data <= 'd1; 9712: data <= 'd1; 9713: data <= 'd1; 9714: data <= 'd1; 9715: data <= 'd3; 9716: data <= 'd2; 9717: data <= 'd0; 9718: data <= 'd0; 9719: data <= 'd0; 9720: data <= 'd0; 9721: data <= 'd0; 9722: data <= 'd0; 9723: data <= 'd0; 9724: data <= 'd0; 9725: data <= 'd0; 9726: data <= 'd0; 9727: data <= 'd0; 9728: data <= 'd0; 9729: data <= 'd0; 9730: data <= 'd0; 9731: data <= 'd0; 9732: data <= 'd0; 9733: data <= 'd2; 9734: data <= 'd5; 9735: data <= 'd3; 9736: data <= 'd1; 9737: data <= 'd1; 9738: data <= 'd1; 9739: data <= 'd5; 9740: data <= 'd5; 9741: data <= 'd5; 9742: data <= 'd5; 9743: data <= 'd5; 9744: data <= 'd5; 9745: data <= 'd5; 9746: data <= 'd1; 9747: data <= 'd1; 9748: data <= 'd2; 9749: data <= 'd0; 9750: data <= 'd0; 9751: data <= 'd0; 9752: data <= 'd0; 9753: data <= 'd0; 9754: data <= 'd0; 9755: data <= 'd0; 9756: data <= 'd0; 9757: data <= 'd0; 9758: data <= 'd0; 9759: data <= 'd0; 9760: data <= 'd0; 9761: data <= 'd0; 9762: data <= 'd0; 9763: data <= 'd0; 9764: data <= 'd0; 9765: data <= 'd2; 9766: data <= 'd6; 9767: data <= 'd1; 9768: data <= 'd5; 9769: data <= 'd2; 9770: data <= 'd2; 9771: data <= 'd2; 9772: data <= 'd2; 9773: data <= 'd2; 9774: data <= 'd2; 9775: data <= 'd2; 9776: data <= 'd2; 9777: data <= 'd2; 9778: data <= 'd2; 9779: data <= 'd5; 9780: data <= 'd2; 9781: data <= 'd0; 9782: data <= 'd0; 9783: data <= 'd0; 9784: data <= 'd0; 9785: data <= 'd0; 9786: data <= 'd0; 9787: data <= 'd0; 9788: data <= 'd0; 9789: data <= 'd0; 9790: data <= 'd0; 9791: data <= 'd0; 9792: data <= 'd0; 9793: data <= 'd0; 9794: data <= 'd0; 9795: data <= 'd2; 9796: data <= 'd2; 9797: data <= 'd2; 9798: data <= 'd1; 9799: data <= 'd5; 9800: data <= 'd2; 9801: data <= 'd8; 9802: data <= 'd8; 9803: data <= 'd8; 9804: data <= 'd8; 9805: data <= 'd8; 9806: data <= 'd9; 9807: data <= 'd9; 9808: data <= 'd8; 9809: data <= 'd8; 9810: data <= 'd8; 9811: data <= 'd2; 9812: data <= 'd2; 9813: data <= 'd0; 9814: data <= 'd0; 9815: data <= 'd0; 9816: data <= 'd0; 9817: data <= 'd0; 9818: data <= 'd0; 9819: data <= 'd0; 9820: data <= 'd0; 9821: data <= 'd0; 9822: data <= 'd0; 9823: data <= 'd0; 9824: data <= 'd0; 9825: data <= 'd0; 9826: data <= 'd0; 9827: data <= 'd2; 9828: data <= 'd1; 9829: data <= 'd2; 9830: data <= 'd1; 9831: data <= 'd2; 9832: data <= 'd8; 9833: data <= 'd8; 9834: data <= 'd9; 9835: data <= 'd9; 9836: data <= 'd2; 9837: data <= 'd9; 9838: data <= 'd11; 9839: data <= 'd11; 9840: data <= 'd10; 9841: data <= 'd2; 9842: data <= 'd9; 9843: data <= 'd2; 9844: data <= 'd2; 9845: data <= 'd0; 9846: data <= 'd0; 9847: data <= 'd0; 9848: data <= 'd0; 9849: data <= 'd0; 9850: data <= 'd0; 9851: data <= 'd0; 9852: data <= 'd0; 9853: data <= 'd0; 9854: data <= 'd0; 9855: data <= 'd0; 9856: data <= 'd0; 9857: data <= 'd0; 9858: data <= 'd0; 9859: data <= 'd2; 9860: data <= 'd5; 9861: data <= 'd1; 9862: data <= 'd2; 9863: data <= 'd9; 9864: data <= 'd10; 9865: data <= 'd9; 9866: data <= 'd9; 9867: data <= 'd10; 9868: data <= 'd11; 9869: data <= 'd10; 9870: data <= 'd11; 9871: data <= 'd11; 9872: data <= 'd10; 9873: data <= 'd11; 9874: data <= 'd10; 9875: data <= 'd9; 9876: data <= 'd2; 9877: data <= 'd0; 9878: data <= 'd0; 9879: data <= 'd0; 9880: data <= 'd0; 9881: data <= 'd0; 9882: data <= 'd0; 9883: data <= 'd0; 9884: data <= 'd0; 9885: data <= 'd0; 9886: data <= 'd0; 9887: data <= 'd0; 9888: data <= 'd0; 9889: data <= 'd0; 9890: data <= 'd0; 9891: data <= 'd0; 9892: data <= 'd2; 9893: data <= 'd5; 9894: data <= 'd5; 9895: data <= 'd2; 9896: data <= 'd8; 9897: data <= 'd9; 9898: data <= 'd9; 9899: data <= 'd10; 9900: data <= 'd10; 9901: data <= 'd10; 9902: data <= 'd8; 9903: data <= 'd8; 9904: data <= 'd10; 9905: data <= 'd10; 9906: data <= 'd9; 9907: data <= 'd2; 9908: data <= 'd0; 9909: data <= 'd0; 9910: data <= 'd0; 9911: data <= 'd0; 9912: data <= 'd0; 9913: data <= 'd0; 9914: data <= 'd0; 9915: data <= 'd0; 9916: data <= 'd0; 9917: data <= 'd0; 9918: data <= 'd0; 9919: data <= 'd0; 9920: data <= 'd0; 9921: data <= 'd0; 9922: data <= 'd0; 9923: data <= 'd0; 9924: data <= 'd0; 9925: data <= 'd2; 9926: data <= 'd2; 9927: data <= 'd2; 9928: data <= 'd5; 9929: data <= 'd8; 9930: data <= 'd9; 9931: data <= 'd9; 9932: data <= 'd10; 9933: data <= 'd10; 9934: data <= 'd9; 9935: data <= 'd9; 9936: data <= 'd10; 9937: data <= 'd10; 9938: data <= 'd9; 9939: data <= 'd2; 9940: data <= 'd0; 9941: data <= 'd0; 9942: data <= 'd0; 9943: data <= 'd0; 9944: data <= 'd0; 9945: data <= 'd0; 9946: data <= 'd0; 9947: data <= 'd0; 9948: data <= 'd0; 9949: data <= 'd0; 9950: data <= 'd0; 9951: data <= 'd0; 9952: data <= 'd0; 9953: data <= 'd0; 9954: data <= 'd0; 9955: data <= 'd0; 9956: data <= 'd0; 9957: data <= 'd0; 9958: data <= 'd0; 9959: data <= 'd0; 9960: data <= 'd2; 9961: data <= 'd5; 9962: data <= 'd5; 9963: data <= 'd8; 9964: data <= 'd9; 9965: data <= 'd9; 9966: data <= 'd9; 9967: data <= 'd9; 9968: data <= 'd9; 9969: data <= 'd9; 9970: data <= 'd5; 9971: data <= 'd2; 9972: data <= 'd0; 9973: data <= 'd0; 9974: data <= 'd0; 9975: data <= 'd0; 9976: data <= 'd0; 9977: data <= 'd0; 9978: data <= 'd0; 9979: data <= 'd0; 9980: data <= 'd0; 9981: data <= 'd0; 9982: data <= 'd0; 9983: data <= 'd0; 9984: data <= 'd0; 9985: data <= 'd0; 9986: data <= 'd0; 9987: data <= 'd0; 9988: data <= 'd0; 9989: data <= 'd0; 9990: data <= 'd0; 9991: data <= 'd2; 9992: data <= 'd7; 9993: data <= 'd1; 9994: data <= 'd1; 9995: data <= 'd3; 9996: data <= 'd3; 9997: data <= 'd3; 9998: data <= 'd5; 9999: data <= 'd5; 10000: data <= 'd3; 10001: data <= 'd3; 10002: data <= 'd1; 10003: data <= 'd2; 10004: data <= 'd2; 10005: data <= 'd2; 10006: data <= 'd0; 10007: data <= 'd0; 10008: data <= 'd0; 10009: data <= 'd0; 10010: data <= 'd0; 10011: data <= 'd0; 10012: data <= 'd0; 10013: data <= 'd0; 10014: data <= 'd0; 10015: data <= 'd0; 10016: data <= 'd0; 10017: data <= 'd0; 10018: data <= 'd0; 10019: data <= 'd0; 10020: data <= 'd0; 10021: data <= 'd0; 10022: data <= 'd0; 10023: data <= 'd2; 10024: data <= 'd7; 10025: data <= 'd7; 10026: data <= 'd5; 10027: data <= 'd3; 10028: data <= 'd3; 10029: data <= 'd3; 10030: data <= 'd1; 10031: data <= 'd1; 10032: data <= 'd3; 10033: data <= 'd3; 10034: data <= 'd1; 10035: data <= 'd4; 10036: data <= 'd9; 10037: data <= 'd9; 10038: data <= 'd2; 10039: data <= 'd0; 10040: data <= 'd0; 10041: data <= 'd0; 10042: data <= 'd0; 10043: data <= 'd0; 10044: data <= 'd0; 10045: data <= 'd0; 10046: data <= 'd0; 10047: data <= 'd0; 10048: data <= 'd0; 10049: data <= 'd0; 10050: data <= 'd0; 10051: data <= 'd0; 10052: data <= 'd0; 10053: data <= 'd0; 10054: data <= 'd0; 10055: data <= 'd2; 10056: data <= 'd4; 10057: data <= 'd9; 10058: data <= 'd9; 10059: data <= 'd1; 10060: data <= 'd3; 10061: data <= 'd3; 10062: data <= 'd1; 10063: data <= 'd1; 10064: data <= 'd3; 10065: data <= 'd1; 10066: data <= 'd1; 10067: data <= 'd4; 10068: data <= 'd9; 10069: data <= 'd9; 10070: data <= 'd2; 10071: data <= 'd0; 10072: data <= 'd0; 10073: data <= 'd0; 10074: data <= 'd0; 10075: data <= 'd0; 10076: data <= 'd0; 10077: data <= 'd0; 10078: data <= 'd0; 10079: data <= 'd0; 10080: data <= 'd0; 10081: data <= 'd0; 10082: data <= 'd0; 10083: data <= 'd0; 10084: data <= 'd0; 10085: data <= 'd0; 10086: data <= 'd0; 10087: data <= 'd0; 10088: data <= 'd2; 10089: data <= 'd9; 10090: data <= 'd9; 10091: data <= 'd2; 10092: data <= 'd2; 10093: data <= 'd5; 10094: data <= 'd5; 10095: data <= 'd5; 10096: data <= 'd2; 10097: data <= 'd2; 10098: data <= 'd2; 10099: data <= 'd5; 10100: data <= 'd2; 10101: data <= 'd2; 10102: data <= 'd0; 10103: data <= 'd0; 10104: data <= 'd0; 10105: data <= 'd0; 10106: data <= 'd0; 10107: data <= 'd0; 10108: data <= 'd0; 10109: data <= 'd0; 10110: data <= 'd0; 10111: data <= 'd0; 10112: data <= 'd0; 10113: data <= 'd0; 10114: data <= 'd0; 10115: data <= 'd0; 10116: data <= 'd0; 10117: data <= 'd0; 10118: data <= 'd0; 10119: data <= 'd0; 10120: data <= 'd2; 10121: data <= 'd2; 10122: data <= 'd2; 10123: data <= 'd1; 10124: data <= 'd3; 10125: data <= 'd3; 10126: data <= 'd1; 10127: data <= 'd3; 10128: data <= 'd3; 10129: data <= 'd3; 10130: data <= 'd2; 10131: data <= 'd2; 10132: data <= 'd0; 10133: data <= 'd0; 10134: data <= 'd0; 10135: data <= 'd0; 10136: data <= 'd0; 10137: data <= 'd0; 10138: data <= 'd0; 10139: data <= 'd0; 10140: data <= 'd0; 10141: data <= 'd0; 10142: data <= 'd0; 10143: data <= 'd0; 10144: data <= 'd0; 10145: data <= 'd0; 10146: data <= 'd0; 10147: data <= 'd0; 10148: data <= 'd0; 10149: data <= 'd0; 10150: data <= 'd0; 10151: data <= 'd0; 10152: data <= 'd2; 10153: data <= 'd4; 10154: data <= 'd7; 10155: data <= 'd7; 10156: data <= 'd2; 10157: data <= 'd2; 10158: data <= 'd2; 10159: data <= 'd5; 10160: data <= 'd5; 10161: data <= 'd4; 10162: data <= 'd2; 10163: data <= 'd0; 10164: data <= 'd0; 10165: data <= 'd0; 10166: data <= 'd0; 10167: data <= 'd0; 10168: data <= 'd0; 10169: data <= 'd0; 10170: data <= 'd0; 10171: data <= 'd0; 10172: data <= 'd0; 10173: data <= 'd0; 10174: data <= 'd0; 10175: data <= 'd0; 10176: data <= 'd0; 10177: data <= 'd0; 10178: data <= 'd0; 10179: data <= 'd0; 10180: data <= 'd0; 10181: data <= 'd0; 10182: data <= 'd0; 10183: data <= 'd0; 10184: data <= 'd0; 10185: data <= 'd2; 10186: data <= 'd4; 10187: data <= 'd7; 10188: data <= 'd2; 10189: data <= 'd0; 10190: data <= 'd0; 10191: data <= 'd2; 10192: data <= 'd4; 10193: data <= 'd4; 10194: data <= 'd2; 10195: data <= 'd0; 10196: data <= 'd0; 10197: data <= 'd0; 10198: data <= 'd0; 10199: data <= 'd0; 10200: data <= 'd0; 10201: data <= 'd0; 10202: data <= 'd0; 10203: data <= 'd0; 10204: data <= 'd0; 10205: data <= 'd0; 10206: data <= 'd0; 10207: data <= 'd0; 10208: data <= 'd0; 10209: data <= 'd0; 10210: data <= 'd0; 10211: data <= 'd0; 10212: data <= 'd0; 10213: data <= 'd0; 10214: data <= 'd0; 10215: data <= 'd0; 10216: data <= 'd0; 10217: data <= 'd2; 10218: data <= 'd2; 10219: data <= 'd2; 10220: data <= 'd2; 10221: data <= 'd0; 10222: data <= 'd0; 10223: data <= 'd0; 10224: data <= 'd2; 10225: data <= 'd2; 10226: data <= 'd2; 10227: data <= 'd0; 10228: data <= 'd0; 10229: data <= 'd0; 10230: data <= 'd0; 10231: data <= 'd0; 10232: data <= 'd0; 10233: data <= 'd0; 10234: data <= 'd0; 10235: data <= 'd0; 10236: data <= 'd0; 10237: data <= 'd0; 10238: data <= 'd0; 10239: data <= 'd0; 10240: data <= 'd0; 10241: data <= 'd0; 10242: data <= 'd0; 10243: data <= 'd0; 10244: data <= 'd0; 10245: data <= 'd0; 10246: data <= 'd0; 10247: data <= 'd0; 10248: data <= 'd0; 10249: data <= 'd0; 10250: data <= 'd0; 10251: data <= 'd0; 10252: data <= 'd0; 10253: data <= 'd0; 10254: data <= 'd0; 10255: data <= 'd0; 10256: data <= 'd0; 10257: data <= 'd0; 10258: data <= 'd0; 10259: data <= 'd0; 10260: data <= 'd0; 10261: data <= 'd0; 10262: data <= 'd0; 10263: data <= 'd0; 10264: data <= 'd0; 10265: data <= 'd0; 10266: data <= 'd0; 10267: data <= 'd0; 10268: data <= 'd0; 10269: data <= 'd0; 10270: data <= 'd0; 10271: data <= 'd0; 10272: data <= 'd0; 10273: data <= 'd0; 10274: data <= 'd0; 10275: data <= 'd0; 10276: data <= 'd0; 10277: data <= 'd0; 10278: data <= 'd0; 10279: data <= 'd0; 10280: data <= 'd0; 10281: data <= 'd0; 10282: data <= 'd0; 10283: data <= 'd0; 10284: data <= 'd0; 10285: data <= 'd0; 10286: data <= 'd0; 10287: data <= 'd0; 10288: data <= 'd0; 10289: data <= 'd0; 10290: data <= 'd0; 10291: data <= 'd0; 10292: data <= 'd0; 10293: data <= 'd0; 10294: data <= 'd0; 10295: data <= 'd0; 10296: data <= 'd0; 10297: data <= 'd0; 10298: data <= 'd0; 10299: data <= 'd0; 10300: data <= 'd0; 10301: data <= 'd0; 10302: data <= 'd0; 10303: data <= 'd0; 10304: data <= 'd0; 10305: data <= 'd0; 10306: data <= 'd0; 10307: data <= 'd0; 10308: data <= 'd0; 10309: data <= 'd0; 10310: data <= 'd0; 10311: data <= 'd0; 10312: data <= 'd0; 10313: data <= 'd0; 10314: data <= 'd0; 10315: data <= 'd0; 10316: data <= 'd0; 10317: data <= 'd0; 10318: data <= 'd0; 10319: data <= 'd0; 10320: data <= 'd0; 10321: data <= 'd0; 10322: data <= 'd0; 10323: data <= 'd0; 10324: data <= 'd0; 10325: data <= 'd0; 10326: data <= 'd0; 10327: data <= 'd0; 10328: data <= 'd0; 10329: data <= 'd0; 10330: data <= 'd0; 10331: data <= 'd0; 10332: data <= 'd0; 10333: data <= 'd0; 10334: data <= 'd0; 10335: data <= 'd0; 10336: data <= 'd0; 10337: data <= 'd0; 10338: data <= 'd0; 10339: data <= 'd0; 10340: data <= 'd0; 10341: data <= 'd0; 10342: data <= 'd0; 10343: data <= 'd0; 10344: data <= 'd0; 10345: data <= 'd0; 10346: data <= 'd0; 10347: data <= 'd0; 10348: data <= 'd0; 10349: data <= 'd0; 10350: data <= 'd0; 10351: data <= 'd0; 10352: data <= 'd0; 10353: data <= 'd0; 10354: data <= 'd0; 10355: data <= 'd0; 10356: data <= 'd0; 10357: data <= 'd0; 10358: data <= 'd0; 10359: data <= 'd0; 10360: data <= 'd0; 10361: data <= 'd0; 10362: data <= 'd0; 10363: data <= 'd0; 10364: data <= 'd0; 10365: data <= 'd0; 10366: data <= 'd0; 10367: data <= 'd0; 10368: data <= 'd0; 10369: data <= 'd0; 10370: data <= 'd0; 10371: data <= 'd0; 10372: data <= 'd0; 10373: data <= 'd0; 10374: data <= 'd0; 10375: data <= 'd0; 10376: data <= 'd0; 10377: data <= 'd0; 10378: data <= 'd0; 10379: data <= 'd0; 10380: data <= 'd0; 10381: data <= 'd0; 10382: data <= 'd0; 10383: data <= 'd0; 10384: data <= 'd0; 10385: data <= 'd0; 10386: data <= 'd0; 10387: data <= 'd0; 10388: data <= 'd0; 10389: data <= 'd0; 10390: data <= 'd0; 10391: data <= 'd0; 10392: data <= 'd0; 10393: data <= 'd0; 10394: data <= 'd0; 10395: data <= 'd0; 10396: data <= 'd0; 10397: data <= 'd0; 10398: data <= 'd0; 10399: data <= 'd0; 10400: data <= 'd0; 10401: data <= 'd0; 10402: data <= 'd0; 10403: data <= 'd0; 10404: data <= 'd0; 10405: data <= 'd0; 10406: data <= 'd0; 10407: data <= 'd0; 10408: data <= 'd0; 10409: data <= 'd0; 10410: data <= 'd0; 10411: data <= 'd0; 10412: data <= 'd0; 10413: data <= 'd0; 10414: data <= 'd0; 10415: data <= 'd0; 10416: data <= 'd0; 10417: data <= 'd0; 10418: data <= 'd0; 10419: data <= 'd0; 10420: data <= 'd0; 10421: data <= 'd0; 10422: data <= 'd0; 10423: data <= 'd0; 10424: data <= 'd0; 10425: data <= 'd0; 10426: data <= 'd0; 10427: data <= 'd0; 10428: data <= 'd0; 10429: data <= 'd0; 10430: data <= 'd0; 10431: data <= 'd0; 10432: data <= 'd0; 10433: data <= 'd0; 10434: data <= 'd0; 10435: data <= 'd0; 10436: data <= 'd0; 10437: data <= 'd0; 10438: data <= 'd0; 10439: data <= 'd0; 10440: data <= 'd0; 10441: data <= 'd0; 10442: data <= 'd0; 10443: data <= 'd0; 10444: data <= 'd0; 10445: data <= 'd0; 10446: data <= 'd0; 10447: data <= 'd0; 10448: data <= 'd0; 10449: data <= 'd0; 10450: data <= 'd0; 10451: data <= 'd0; 10452: data <= 'd0; 10453: data <= 'd0; 10454: data <= 'd0; 10455: data <= 'd0; 10456: data <= 'd0; 10457: data <= 'd0; 10458: data <= 'd0; 10459: data <= 'd0; 10460: data <= 'd0; 10461: data <= 'd0; 10462: data <= 'd0; 10463: data <= 'd0; 10464: data <= 'd0; 10465: data <= 'd0; 10466: data <= 'd0; 10467: data <= 'd0; 10468: data <= 'd0; 10469: data <= 'd0; 10470: data <= 'd0; 10471: data <= 'd0; 10472: data <= 'd0; 10473: data <= 'd0; 10474: data <= 'd0; 10475: data <= 'd0; 10476: data <= 'd0; 10477: data <= 'd0; 10478: data <= 'd0; 10479: data <= 'd0; 10480: data <= 'd0; 10481: data <= 'd0; 10482: data <= 'd0; 10483: data <= 'd0; 10484: data <= 'd0; 10485: data <= 'd0; 10486: data <= 'd0; 10487: data <= 'd0; 10488: data <= 'd0; 10489: data <= 'd0; 10490: data <= 'd0; 10491: data <= 'd0; 10492: data <= 'd0; 10493: data <= 'd0; 10494: data <= 'd0; 10495: data <= 'd0; 10496: data <= 'd0; 10497: data <= 'd0; 10498: data <= 'd0; 10499: data <= 'd0; 10500: data <= 'd0; 10501: data <= 'd0; 10502: data <= 'd0; 10503: data <= 'd0; 10504: data <= 'd0; 10505: data <= 'd0; 10506: data <= 'd0; 10507: data <= 'd0; 10508: data <= 'd0; 10509: data <= 'd0; 10510: data <= 'd0; 10511: data <= 'd0; 10512: data <= 'd0; 10513: data <= 'd0; 10514: data <= 'd0; 10515: data <= 'd0; 10516: data <= 'd0; 10517: data <= 'd0; 10518: data <= 'd0; 10519: data <= 'd0; 10520: data <= 'd0; 10521: data <= 'd0; 10522: data <= 'd0; 10523: data <= 'd0; 10524: data <= 'd0; 10525: data <= 'd0; 10526: data <= 'd0; 10527: data <= 'd0; 10528: data <= 'd0; 10529: data <= 'd0; 10530: data <= 'd0; 10531: data <= 'd0; 10532: data <= 'd0; 10533: data <= 'd0; 10534: data <= 'd0; 10535: data <= 'd0; 10536: data <= 'd0; 10537: data <= 'd0; 10538: data <= 'd0; 10539: data <= 'd0; 10540: data <= 'd0; 10541: data <= 'd2; 10542: data <= 'd2; 10543: data <= 'd2; 10544: data <= 'd2; 10545: data <= 'd2; 10546: data <= 'd2; 10547: data <= 'd0; 10548: data <= 'd0; 10549: data <= 'd0; 10550: data <= 'd0; 10551: data <= 'd0; 10552: data <= 'd0; 10553: data <= 'd0; 10554: data <= 'd0; 10555: data <= 'd0; 10556: data <= 'd0; 10557: data <= 'd0; 10558: data <= 'd0; 10559: data <= 'd0; 10560: data <= 'd0; 10561: data <= 'd0; 10562: data <= 'd0; 10563: data <= 'd0; 10564: data <= 'd0; 10565: data <= 'd0; 10566: data <= 'd0; 10567: data <= 'd0; 10568: data <= 'd0; 10569: data <= 'd0; 10570: data <= 'd0; 10571: data <= 'd2; 10572: data <= 'd2; 10573: data <= 'd6; 10574: data <= 'd6; 10575: data <= 'd6; 10576: data <= 'd6; 10577: data <= 'd6; 10578: data <= 'd6; 10579: data <= 'd2; 10580: data <= 'd2; 10581: data <= 'd0; 10582: data <= 'd0; 10583: data <= 'd0; 10584: data <= 'd0; 10585: data <= 'd0; 10586: data <= 'd0; 10587: data <= 'd0; 10588: data <= 'd0; 10589: data <= 'd0; 10590: data <= 'd0; 10591: data <= 'd0; 10592: data <= 'd0; 10593: data <= 'd0; 10594: data <= 'd0; 10595: data <= 'd0; 10596: data <= 'd0; 10597: data <= 'd0; 10598: data <= 'd0; 10599: data <= 'd0; 10600: data <= 'd0; 10601: data <= 'd0; 10602: data <= 'd2; 10603: data <= 'd1; 10604: data <= 'd3; 10605: data <= 'd6; 10606: data <= 'd6; 10607: data <= 'd6; 10608: data <= 'd6; 10609: data <= 'd6; 10610: data <= 'd6; 10611: data <= 'd6; 10612: data <= 'd3; 10613: data <= 'd2; 10614: data <= 'd0; 10615: data <= 'd0; 10616: data <= 'd0; 10617: data <= 'd0; 10618: data <= 'd0; 10619: data <= 'd0; 10620: data <= 'd0; 10621: data <= 'd0; 10622: data <= 'd0; 10623: data <= 'd0; 10624: data <= 'd0; 10625: data <= 'd0; 10626: data <= 'd0; 10627: data <= 'd0; 10628: data <= 'd0; 10629: data <= 'd0; 10630: data <= 'd0; 10631: data <= 'd0; 10632: data <= 'd0; 10633: data <= 'd2; 10634: data <= 'd1; 10635: data <= 'd1; 10636: data <= 'd1; 10637: data <= 'd3; 10638: data <= 'd6; 10639: data <= 'd6; 10640: data <= 'd6; 10641: data <= 'd6; 10642: data <= 'd6; 10643: data <= 'd3; 10644: data <= 'd1; 10645: data <= 'd1; 10646: data <= 'd2; 10647: data <= 'd0; 10648: data <= 'd0; 10649: data <= 'd0; 10650: data <= 'd0; 10651: data <= 'd0; 10652: data <= 'd0; 10653: data <= 'd0; 10654: data <= 'd0; 10655: data <= 'd0; 10656: data <= 'd0; 10657: data <= 'd0; 10658: data <= 'd0; 10659: data <= 'd0; 10660: data <= 'd0; 10661: data <= 'd0; 10662: data <= 'd0; 10663: data <= 'd0; 10664: data <= 'd0; 10665: data <= 'd2; 10666: data <= 'd1; 10667: data <= 'd1; 10668: data <= 'd5; 10669: data <= 'd5; 10670: data <= 'd5; 10671: data <= 'd1; 10672: data <= 'd1; 10673: data <= 'd1; 10674: data <= 'd1; 10675: data <= 'd1; 10676: data <= 'd5; 10677: data <= 'd5; 10678: data <= 'd2; 10679: data <= 'd0; 10680: data <= 'd0; 10681: data <= 'd0; 10682: data <= 'd0; 10683: data <= 'd0; 10684: data <= 'd0; 10685: data <= 'd0; 10686: data <= 'd0; 10687: data <= 'd0; 10688: data <= 'd0; 10689: data <= 'd0; 10690: data <= 'd0; 10691: data <= 'd0; 10692: data <= 'd0; 10693: data <= 'd0; 10694: data <= 'd0; 10695: data <= 'd0; 10696: data <= 'd2; 10697: data <= 'd1; 10698: data <= 'd5; 10699: data <= 'd5; 10700: data <= 'd3; 10701: data <= 'd6; 10702: data <= 'd6; 10703: data <= 'd6; 10704: data <= 'd6; 10705: data <= 'd6; 10706: data <= 'd6; 10707: data <= 'd6; 10708: data <= 'd6; 10709: data <= 'd3; 10710: data <= 'd5; 10711: data <= 'd2; 10712: data <= 'd0; 10713: data <= 'd0; 10714: data <= 'd0; 10715: data <= 'd0; 10716: data <= 'd0; 10717: data <= 'd0; 10718: data <= 'd0; 10719: data <= 'd0; 10720: data <= 'd0; 10721: data <= 'd0; 10722: data <= 'd0; 10723: data <= 'd0; 10724: data <= 'd0; 10725: data <= 'd0; 10726: data <= 'd0; 10727: data <= 'd0; 10728: data <= 'd2; 10729: data <= 'd5; 10730: data <= 'd3; 10731: data <= 'd6; 10732: data <= 'd3; 10733: data <= 'd1; 10734: data <= 'd1; 10735: data <= 'd1; 10736: data <= 'd1; 10737: data <= 'd1; 10738: data <= 'd1; 10739: data <= 'd1; 10740: data <= 'd1; 10741: data <= 'd1; 10742: data <= 'd3; 10743: data <= 'd2; 10744: data <= 'd0; 10745: data <= 'd0; 10746: data <= 'd0; 10747: data <= 'd0; 10748: data <= 'd0; 10749: data <= 'd0; 10750: data <= 'd0; 10751: data <= 'd0; 10752: data <= 'd0; 10753: data <= 'd0; 10754: data <= 'd0; 10755: data <= 'd0; 10756: data <= 'd0; 10757: data <= 'd0; 10758: data <= 'd0; 10759: data <= 'd0; 10760: data <= 'd2; 10761: data <= 'd5; 10762: data <= 'd3; 10763: data <= 'd1; 10764: data <= 'd1; 10765: data <= 'd1; 10766: data <= 'd5; 10767: data <= 'd5; 10768: data <= 'd5; 10769: data <= 'd5; 10770: data <= 'd5; 10771: data <= 'd5; 10772: data <= 'd5; 10773: data <= 'd1; 10774: data <= 'd1; 10775: data <= 'd2; 10776: data <= 'd0; 10777: data <= 'd0; 10778: data <= 'd0; 10779: data <= 'd0; 10780: data <= 'd0; 10781: data <= 'd0; 10782: data <= 'd0; 10783: data <= 'd0; 10784: data <= 'd0; 10785: data <= 'd0; 10786: data <= 'd0; 10787: data <= 'd0; 10788: data <= 'd0; 10789: data <= 'd0; 10790: data <= 'd0; 10791: data <= 'd0; 10792: data <= 'd2; 10793: data <= 'd6; 10794: data <= 'd1; 10795: data <= 'd5; 10796: data <= 'd2; 10797: data <= 'd2; 10798: data <= 'd2; 10799: data <= 'd2; 10800: data <= 'd2; 10801: data <= 'd2; 10802: data <= 'd2; 10803: data <= 'd2; 10804: data <= 'd2; 10805: data <= 'd2; 10806: data <= 'd5; 10807: data <= 'd2; 10808: data <= 'd0; 10809: data <= 'd0; 10810: data <= 'd0; 10811: data <= 'd0; 10812: data <= 'd0; 10813: data <= 'd0; 10814: data <= 'd0; 10815: data <= 'd0; 10816: data <= 'd0; 10817: data <= 'd0; 10818: data <= 'd0; 10819: data <= 'd0; 10820: data <= 'd0; 10821: data <= 'd0; 10822: data <= 'd2; 10823: data <= 'd2; 10824: data <= 'd2; 10825: data <= 'd1; 10826: data <= 'd5; 10827: data <= 'd2; 10828: data <= 'd8; 10829: data <= 'd8; 10830: data <= 'd8; 10831: data <= 'd8; 10832: data <= 'd8; 10833: data <= 'd9; 10834: data <= 'd9; 10835: data <= 'd8; 10836: data <= 'd8; 10837: data <= 'd8; 10838: data <= 'd2; 10839: data <= 'd2; 10840: data <= 'd0; 10841: data <= 'd0; 10842: data <= 'd0; 10843: data <= 'd0; 10844: data <= 'd0; 10845: data <= 'd0; 10846: data <= 'd0; 10847: data <= 'd0; 10848: data <= 'd0; 10849: data <= 'd0; 10850: data <= 'd0; 10851: data <= 'd0; 10852: data <= 'd0; 10853: data <= 'd0; 10854: data <= 'd2; 10855: data <= 'd1; 10856: data <= 'd2; 10857: data <= 'd1; 10858: data <= 'd2; 10859: data <= 'd8; 10860: data <= 'd8; 10861: data <= 'd9; 10862: data <= 'd9; 10863: data <= 'd2; 10864: data <= 'd9; 10865: data <= 'd11; 10866: data <= 'd11; 10867: data <= 'd10; 10868: data <= 'd2; 10869: data <= 'd9; 10870: data <= 'd2; 10871: data <= 'd2; 10872: data <= 'd0; 10873: data <= 'd0; 10874: data <= 'd0; 10875: data <= 'd0; 10876: data <= 'd0; 10877: data <= 'd0; 10878: data <= 'd0; 10879: data <= 'd0; 10880: data <= 'd0; 10881: data <= 'd0; 10882: data <= 'd0; 10883: data <= 'd0; 10884: data <= 'd0; 10885: data <= 'd0; 10886: data <= 'd2; 10887: data <= 'd5; 10888: data <= 'd1; 10889: data <= 'd2; 10890: data <= 'd9; 10891: data <= 'd10; 10892: data <= 'd9; 10893: data <= 'd9; 10894: data <= 'd10; 10895: data <= 'd11; 10896: data <= 'd10; 10897: data <= 'd11; 10898: data <= 'd11; 10899: data <= 'd10; 10900: data <= 'd11; 10901: data <= 'd10; 10902: data <= 'd9; 10903: data <= 'd2; 10904: data <= 'd0; 10905: data <= 'd0; 10906: data <= 'd0; 10907: data <= 'd0; 10908: data <= 'd0; 10909: data <= 'd0; 10910: data <= 'd0; 10911: data <= 'd0; 10912: data <= 'd0; 10913: data <= 'd0; 10914: data <= 'd0; 10915: data <= 'd0; 10916: data <= 'd0; 10917: data <= 'd0; 10918: data <= 'd0; 10919: data <= 'd2; 10920: data <= 'd5; 10921: data <= 'd5; 10922: data <= 'd2; 10923: data <= 'd8; 10924: data <= 'd9; 10925: data <= 'd2; 10926: data <= 'd2; 10927: data <= 'd10; 10928: data <= 'd10; 10929: data <= 'd8; 10930: data <= 'd8; 10931: data <= 'd10; 10932: data <= 'd10; 10933: data <= 'd9; 10934: data <= 'd2; 10935: data <= 'd0; 10936: data <= 'd0; 10937: data <= 'd0; 10938: data <= 'd0; 10939: data <= 'd0; 10940: data <= 'd0; 10941: data <= 'd0; 10942: data <= 'd0; 10943: data <= 'd0; 10944: data <= 'd0; 10945: data <= 'd0; 10946: data <= 'd0; 10947: data <= 'd0; 10948: data <= 'd0; 10949: data <= 'd0; 10950: data <= 'd0; 10951: data <= 'd0; 10952: data <= 'd2; 10953: data <= 'd2; 10954: data <= 'd2; 10955: data <= 'd8; 10956: data <= 'd2; 10957: data <= 'd9; 10958: data <= 'd9; 10959: data <= 'd2; 10960: data <= 'd10; 10961: data <= 'd9; 10962: data <= 'd9; 10963: data <= 'd10; 10964: data <= 'd10; 10965: data <= 'd9; 10966: data <= 'd2; 10967: data <= 'd0; 10968: data <= 'd0; 10969: data <= 'd0; 10970: data <= 'd0; 10971: data <= 'd0; 10972: data <= 'd0; 10973: data <= 'd0; 10974: data <= 'd0; 10975: data <= 'd0; 10976: data <= 'd0; 10977: data <= 'd0; 10978: data <= 'd0; 10979: data <= 'd0; 10980: data <= 'd0; 10981: data <= 'd0; 10982: data <= 'd0; 10983: data <= 'd0; 10984: data <= 'd0; 10985: data <= 'd0; 10986: data <= 'd2; 10987: data <= 'd2; 10988: data <= 'd1; 10989: data <= 'd9; 10990: data <= 'd9; 10991: data <= 'd2; 10992: data <= 'd9; 10993: data <= 'd9; 10994: data <= 'd9; 10995: data <= 'd9; 10996: data <= 'd9; 10997: data <= 'd5; 10998: data <= 'd2; 10999: data <= 'd0; 11000: data <= 'd0; 11001: data <= 'd0; 11002: data <= 'd0; 11003: data <= 'd0; 11004: data <= 'd0; 11005: data <= 'd0; 11006: data <= 'd0; 11007: data <= 'd0; 11008: data <= 'd0; 11009: data <= 'd0; 11010: data <= 'd0; 11011: data <= 'd0; 11012: data <= 'd0; 11013: data <= 'd0; 11014: data <= 'd0; 11015: data <= 'd0; 11016: data <= 'd0; 11017: data <= 'd0; 11018: data <= 'd2; 11019: data <= 'd1; 11020: data <= 'd1; 11021: data <= 'd1; 11022: data <= 'd2; 11023: data <= 'd3; 11024: data <= 'd3; 11025: data <= 'd5; 11026: data <= 'd5; 11027: data <= 'd3; 11028: data <= 'd3; 11029: data <= 'd1; 11030: data <= 'd2; 11031: data <= 'd0; 11032: data <= 'd0; 11033: data <= 'd0; 11034: data <= 'd0; 11035: data <= 'd0; 11036: data <= 'd0; 11037: data <= 'd0; 11038: data <= 'd0; 11039: data <= 'd0; 11040: data <= 'd0; 11041: data <= 'd0; 11042: data <= 'd0; 11043: data <= 'd0; 11044: data <= 'd0; 11045: data <= 'd0; 11046: data <= 'd0; 11047: data <= 'd0; 11048: data <= 'd0; 11049: data <= 'd0; 11050: data <= 'd2; 11051: data <= 'd1; 11052: data <= 'd1; 11053: data <= 'd1; 11054: data <= 'd3; 11055: data <= 'd3; 11056: data <= 'd3; 11057: data <= 'd1; 11058: data <= 'd1; 11059: data <= 'd3; 11060: data <= 'd3; 11061: data <= 'd1; 11062: data <= 'd2; 11063: data <= 'd0; 11064: data <= 'd0; 11065: data <= 'd0; 11066: data <= 'd0; 11067: data <= 'd0; 11068: data <= 'd0; 11069: data <= 'd0; 11070: data <= 'd0; 11071: data <= 'd0; 11072: data <= 'd0; 11073: data <= 'd0; 11074: data <= 'd0; 11075: data <= 'd0; 11076: data <= 'd0; 11077: data <= 'd0; 11078: data <= 'd0; 11079: data <= 'd0; 11080: data <= 'd0; 11081: data <= 'd0; 11082: data <= 'd2; 11083: data <= 'd2; 11084: data <= 'd1; 11085: data <= 'd1; 11086: data <= 'd1; 11087: data <= 'd3; 11088: data <= 'd3; 11089: data <= 'd1; 11090: data <= 'd1; 11091: data <= 'd3; 11092: data <= 'd1; 11093: data <= 'd1; 11094: data <= 'd2; 11095: data <= 'd0; 11096: data <= 'd0; 11097: data <= 'd0; 11098: data <= 'd0; 11099: data <= 'd0; 11100: data <= 'd0; 11101: data <= 'd0; 11102: data <= 'd0; 11103: data <= 'd0; 11104: data <= 'd0; 11105: data <= 'd0; 11106: data <= 'd0; 11107: data <= 'd0; 11108: data <= 'd0; 11109: data <= 'd0; 11110: data <= 'd0; 11111: data <= 'd0; 11112: data <= 'd0; 11113: data <= 'd0; 11114: data <= 'd2; 11115: data <= 'd2; 11116: data <= 'd2; 11117: data <= 'd2; 11118: data <= 'd2; 11119: data <= 'd2; 11120: data <= 'd5; 11121: data <= 'd5; 11122: data <= 'd5; 11123: data <= 'd2; 11124: data <= 'd2; 11125: data <= 'd2; 11126: data <= 'd2; 11127: data <= 'd0; 11128: data <= 'd0; 11129: data <= 'd0; 11130: data <= 'd0; 11131: data <= 'd0; 11132: data <= 'd0; 11133: data <= 'd0; 11134: data <= 'd0; 11135: data <= 'd0; 11136: data <= 'd0; 11137: data <= 'd0; 11138: data <= 'd0; 11139: data <= 'd0; 11140: data <= 'd0; 11141: data <= 'd0; 11142: data <= 'd0; 11143: data <= 'd0; 11144: data <= 'd0; 11145: data <= 'd0; 11146: data <= 'd0; 11147: data <= 'd2; 11148: data <= 'd1; 11149: data <= 'd1; 11150: data <= 'd3; 11151: data <= 'd3; 11152: data <= 'd3; 11153: data <= 'd1; 11154: data <= 'd3; 11155: data <= 'd3; 11156: data <= 'd3; 11157: data <= 'd2; 11158: data <= 'd0; 11159: data <= 'd0; 11160: data <= 'd0; 11161: data <= 'd0; 11162: data <= 'd0; 11163: data <= 'd0; 11164: data <= 'd0; 11165: data <= 'd0; 11166: data <= 'd0; 11167: data <= 'd0; 11168: data <= 'd0; 11169: data <= 'd0; 11170: data <= 'd0; 11171: data <= 'd0; 11172: data <= 'd0; 11173: data <= 'd0; 11174: data <= 'd0; 11175: data <= 'd0; 11176: data <= 'd0; 11177: data <= 'd0; 11178: data <= 'd0; 11179: data <= 'd2; 11180: data <= 'd4; 11181: data <= 'd7; 11182: data <= 'd7; 11183: data <= 'd2; 11184: data <= 'd2; 11185: data <= 'd2; 11186: data <= 'd5; 11187: data <= 'd5; 11188: data <= 'd4; 11189: data <= 'd2; 11190: data <= 'd0; 11191: data <= 'd0; 11192: data <= 'd0; 11193: data <= 'd0; 11194: data <= 'd0; 11195: data <= 'd0; 11196: data <= 'd0; 11197: data <= 'd0; 11198: data <= 'd0; 11199: data <= 'd0; 11200: data <= 'd0; 11201: data <= 'd0; 11202: data <= 'd0; 11203: data <= 'd0; 11204: data <= 'd0; 11205: data <= 'd0; 11206: data <= 'd0; 11207: data <= 'd0; 11208: data <= 'd0; 11209: data <= 'd0; 11210: data <= 'd0; 11211: data <= 'd2; 11212: data <= 'd4; 11213: data <= 'd7; 11214: data <= 'd2; 11215: data <= 'd0; 11216: data <= 'd0; 11217: data <= 'd0; 11218: data <= 'd2; 11219: data <= 'd4; 11220: data <= 'd4; 11221: data <= 'd2; 11222: data <= 'd0; 11223: data <= 'd0; 11224: data <= 'd0; 11225: data <= 'd0; 11226: data <= 'd0; 11227: data <= 'd0; 11228: data <= 'd0; 11229: data <= 'd0; 11230: data <= 'd0; 11231: data <= 'd0; 11232: data <= 'd0; 11233: data <= 'd0; 11234: data <= 'd0; 11235: data <= 'd0; 11236: data <= 'd0; 11237: data <= 'd0; 11238: data <= 'd0; 11239: data <= 'd0; 11240: data <= 'd0; 11241: data <= 'd0; 11242: data <= 'd0; 11243: data <= 'd2; 11244: data <= 'd2; 11245: data <= 'd2; 11246: data <= 'd0; 11247: data <= 'd0; 11248: data <= 'd0; 11249: data <= 'd0; 11250: data <= 'd2; 11251: data <= 'd2; 11252: data <= 'd2; 11253: data <= 'd0; 11254: data <= 'd0; 11255: data <= 'd0; 11256: data <= 'd0; 11257: data <= 'd0; 11258: data <= 'd0; 11259: data <= 'd0; 11260: data <= 'd0; 11261: data <= 'd0; 11262: data <= 'd0; 11263: data <= 'd0; 11264: data <= 'd0; 11265: data <= 'd0; 11266: data <= 'd0; 11267: data <= 'd0; 11268: data <= 'd0; 11269: data <= 'd0; 11270: data <= 'd0; 11271: data <= 'd0; 11272: data <= 'd0; 11273: data <= 'd0; 11274: data <= 'd0; 11275: data <= 'd0; 11276: data <= 'd0; 11277: data <= 'd0; 11278: data <= 'd0; 11279: data <= 'd0; 11280: data <= 'd0; 11281: data <= 'd0; 11282: data <= 'd0; 11283: data <= 'd0; 11284: data <= 'd0; 11285: data <= 'd0; 11286: data <= 'd0; 11287: data <= 'd0; 11288: data <= 'd0; 11289: data <= 'd0; 11290: data <= 'd0; 11291: data <= 'd0; 11292: data <= 'd0; 11293: data <= 'd0; 11294: data <= 'd0; 11295: data <= 'd0; 11296: data <= 'd0; 11297: data <= 'd0; 11298: data <= 'd0; 11299: data <= 'd0; 11300: data <= 'd0; 11301: data <= 'd0; 11302: data <= 'd0; 11303: data <= 'd0; 11304: data <= 'd0; 11305: data <= 'd0; 11306: data <= 'd0; 11307: data <= 'd0; 11308: data <= 'd0; 11309: data <= 'd0; 11310: data <= 'd0; 11311: data <= 'd0; 11312: data <= 'd0; 11313: data <= 'd0; 11314: data <= 'd0; 11315: data <= 'd0; 11316: data <= 'd0; 11317: data <= 'd0; 11318: data <= 'd0; 11319: data <= 'd0; 11320: data <= 'd0; 11321: data <= 'd0; 11322: data <= 'd0; 11323: data <= 'd0; 11324: data <= 'd0; 11325: data <= 'd0; 11326: data <= 'd0; 11327: data <= 'd0; 11328: data <= 'd0; 11329: data <= 'd0; 11330: data <= 'd0; 11331: data <= 'd0; 11332: data <= 'd0; 11333: data <= 'd0; 11334: data <= 'd0; 11335: data <= 'd0; 11336: data <= 'd0; 11337: data <= 'd0; 11338: data <= 'd0; 11339: data <= 'd0; 11340: data <= 'd0; 11341: data <= 'd0; 11342: data <= 'd0; 11343: data <= 'd0; 11344: data <= 'd0; 11345: data <= 'd0; 11346: data <= 'd0; 11347: data <= 'd0; 11348: data <= 'd0; 11349: data <= 'd0; 11350: data <= 'd0; 11351: data <= 'd0; 11352: data <= 'd0; 11353: data <= 'd0; 11354: data <= 'd0; 11355: data <= 'd0; 11356: data <= 'd0; 11357: data <= 'd0; 11358: data <= 'd0; 11359: data <= 'd0; 11360: data <= 'd0; 11361: data <= 'd0; 11362: data <= 'd0; 11363: data <= 'd0; 11364: data <= 'd0; 11365: data <= 'd0; 11366: data <= 'd0; 11367: data <= 'd0; 11368: data <= 'd0; 11369: data <= 'd0; 11370: data <= 'd0; 11371: data <= 'd0; 11372: data <= 'd0; 11373: data <= 'd0; 11374: data <= 'd0; 11375: data <= 'd0; 11376: data <= 'd0; 11377: data <= 'd0; 11378: data <= 'd0; 11379: data <= 'd0; 11380: data <= 'd0; 11381: data <= 'd0; 11382: data <= 'd0; 11383: data <= 'd0; 11384: data <= 'd0; 11385: data <= 'd0; 11386: data <= 'd0; 11387: data <= 'd0; 11388: data <= 'd0; 11389: data <= 'd0; 11390: data <= 'd0; 11391: data <= 'd0; 11392: data <= 'd0; 11393: data <= 'd0; 11394: data <= 'd0; 11395: data <= 'd0; 11396: data <= 'd0; 11397: data <= 'd0; 11398: data <= 'd0; 11399: data <= 'd0; 11400: data <= 'd0; 11401: data <= 'd0; 11402: data <= 'd0; 11403: data <= 'd0; 11404: data <= 'd0; 11405: data <= 'd0; 11406: data <= 'd0; 11407: data <= 'd0; 11408: data <= 'd0; 11409: data <= 'd0; 11410: data <= 'd0; 11411: data <= 'd0; 11412: data <= 'd0; 11413: data <= 'd0; 11414: data <= 'd0; 11415: data <= 'd0; 11416: data <= 'd0; 11417: data <= 'd0; 11418: data <= 'd0; 11419: data <= 'd0; 11420: data <= 'd0; 11421: data <= 'd0; 11422: data <= 'd0; 11423: data <= 'd0; 11424: data <= 'd0; 11425: data <= 'd0; 11426: data <= 'd0; 11427: data <= 'd0; 11428: data <= 'd0; 11429: data <= 'd0; 11430: data <= 'd0; 11431: data <= 'd0; 11432: data <= 'd0; 11433: data <= 'd0; 11434: data <= 'd0; 11435: data <= 'd0; 11436: data <= 'd0; 11437: data <= 'd0; 11438: data <= 'd0; 11439: data <= 'd0; 11440: data <= 'd0; 11441: data <= 'd0; 11442: data <= 'd0; 11443: data <= 'd0; 11444: data <= 'd0; 11445: data <= 'd0; 11446: data <= 'd0; 11447: data <= 'd0; 11448: data <= 'd0; 11449: data <= 'd0; 11450: data <= 'd0; 11451: data <= 'd0; 11452: data <= 'd0; 11453: data <= 'd0; 11454: data <= 'd0; 11455: data <= 'd0; 11456: data <= 'd0; 11457: data <= 'd0; 11458: data <= 'd0; 11459: data <= 'd0; 11460: data <= 'd0; 11461: data <= 'd0; 11462: data <= 'd0; 11463: data <= 'd0; 11464: data <= 'd0; 11465: data <= 'd0; 11466: data <= 'd0; 11467: data <= 'd0; 11468: data <= 'd0; 11469: data <= 'd0; 11470: data <= 'd0; 11471: data <= 'd0; 11472: data <= 'd0; 11473: data <= 'd0; 11474: data <= 'd0; 11475: data <= 'd0; 11476: data <= 'd0; 11477: data <= 'd0; 11478: data <= 'd0; 11479: data <= 'd0; 11480: data <= 'd0; 11481: data <= 'd0; 11482: data <= 'd0; 11483: data <= 'd0; 11484: data <= 'd0; 11485: data <= 'd0; 11486: data <= 'd0; 11487: data <= 'd0; 11488: data <= 'd0; 11489: data <= 'd0; 11490: data <= 'd0; 11491: data <= 'd0; 11492: data <= 'd0; 11493: data <= 'd0; 11494: data <= 'd0; 11495: data <= 'd0; 11496: data <= 'd0; 11497: data <= 'd0; 11498: data <= 'd0; 11499: data <= 'd0; 11500: data <= 'd0; 11501: data <= 'd0; 11502: data <= 'd0; 11503: data <= 'd0; 11504: data <= 'd0; 11505: data <= 'd0; 11506: data <= 'd0; 11507: data <= 'd0; 11508: data <= 'd0; 11509: data <= 'd0; 11510: data <= 'd0; 11511: data <= 'd0; 11512: data <= 'd0; 11513: data <= 'd0; 11514: data <= 'd0; 11515: data <= 'd0; 11516: data <= 'd0; 11517: data <= 'd0; 11518: data <= 'd0; 11519: data <= 'd0; 11520: data <= 'd0; 11521: data <= 'd0; 11522: data <= 'd0; 11523: data <= 'd0; 11524: data <= 'd0; 11525: data <= 'd0; 11526: data <= 'd0; 11527: data <= 'd0; 11528: data <= 'd0; 11529: data <= 'd0; 11530: data <= 'd0; 11531: data <= 'd0; 11532: data <= 'd0; 11533: data <= 'd0; 11534: data <= 'd0; 11535: data <= 'd0; 11536: data <= 'd0; 11537: data <= 'd0; 11538: data <= 'd0; 11539: data <= 'd0; 11540: data <= 'd0; 11541: data <= 'd0; 11542: data <= 'd0; 11543: data <= 'd0; 11544: data <= 'd0; 11545: data <= 'd0; 11546: data <= 'd0; 11547: data <= 'd0; 11548: data <= 'd0; 11549: data <= 'd0; 11550: data <= 'd0; 11551: data <= 'd0; 11552: data <= 'd0; 11553: data <= 'd0; 11554: data <= 'd0; 11555: data <= 'd0; 11556: data <= 'd0; 11557: data <= 'd0; 11558: data <= 'd0; 11559: data <= 'd0; 11560: data <= 'd0; 11561: data <= 'd0; 11562: data <= 'd0; 11563: data <= 'd0; 11564: data <= 'd0; 11565: data <= 'd2; 11566: data <= 'd2; 11567: data <= 'd2; 11568: data <= 'd2; 11569: data <= 'd2; 11570: data <= 'd2; 11571: data <= 'd0; 11572: data <= 'd0; 11573: data <= 'd0; 11574: data <= 'd0; 11575: data <= 'd0; 11576: data <= 'd0; 11577: data <= 'd0; 11578: data <= 'd0; 11579: data <= 'd0; 11580: data <= 'd0; 11581: data <= 'd0; 11582: data <= 'd0; 11583: data <= 'd0; 11584: data <= 'd0; 11585: data <= 'd0; 11586: data <= 'd0; 11587: data <= 'd0; 11588: data <= 'd0; 11589: data <= 'd0; 11590: data <= 'd0; 11591: data <= 'd0; 11592: data <= 'd0; 11593: data <= 'd0; 11594: data <= 'd0; 11595: data <= 'd2; 11596: data <= 'd2; 11597: data <= 'd6; 11598: data <= 'd6; 11599: data <= 'd6; 11600: data <= 'd6; 11601: data <= 'd6; 11602: data <= 'd6; 11603: data <= 'd2; 11604: data <= 'd2; 11605: data <= 'd0; 11606: data <= 'd0; 11607: data <= 'd0; 11608: data <= 'd0; 11609: data <= 'd0; 11610: data <= 'd0; 11611: data <= 'd0; 11612: data <= 'd0; 11613: data <= 'd0; 11614: data <= 'd0; 11615: data <= 'd0; 11616: data <= 'd0; 11617: data <= 'd0; 11618: data <= 'd0; 11619: data <= 'd0; 11620: data <= 'd0; 11621: data <= 'd0; 11622: data <= 'd0; 11623: data <= 'd0; 11624: data <= 'd0; 11625: data <= 'd0; 11626: data <= 'd2; 11627: data <= 'd1; 11628: data <= 'd3; 11629: data <= 'd6; 11630: data <= 'd6; 11631: data <= 'd6; 11632: data <= 'd6; 11633: data <= 'd6; 11634: data <= 'd6; 11635: data <= 'd6; 11636: data <= 'd3; 11637: data <= 'd2; 11638: data <= 'd0; 11639: data <= 'd0; 11640: data <= 'd0; 11641: data <= 'd0; 11642: data <= 'd0; 11643: data <= 'd0; 11644: data <= 'd0; 11645: data <= 'd0; 11646: data <= 'd0; 11647: data <= 'd0; 11648: data <= 'd0; 11649: data <= 'd0; 11650: data <= 'd0; 11651: data <= 'd0; 11652: data <= 'd0; 11653: data <= 'd0; 11654: data <= 'd0; 11655: data <= 'd0; 11656: data <= 'd0; 11657: data <= 'd2; 11658: data <= 'd1; 11659: data <= 'd1; 11660: data <= 'd1; 11661: data <= 'd3; 11662: data <= 'd6; 11663: data <= 'd6; 11664: data <= 'd6; 11665: data <= 'd6; 11666: data <= 'd6; 11667: data <= 'd3; 11668: data <= 'd1; 11669: data <= 'd1; 11670: data <= 'd2; 11671: data <= 'd0; 11672: data <= 'd0; 11673: data <= 'd0; 11674: data <= 'd0; 11675: data <= 'd0; 11676: data <= 'd0; 11677: data <= 'd0; 11678: data <= 'd0; 11679: data <= 'd0; 11680: data <= 'd0; 11681: data <= 'd0; 11682: data <= 'd0; 11683: data <= 'd0; 11684: data <= 'd0; 11685: data <= 'd0; 11686: data <= 'd0; 11687: data <= 'd0; 11688: data <= 'd0; 11689: data <= 'd2; 11690: data <= 'd1; 11691: data <= 'd1; 11692: data <= 'd5; 11693: data <= 'd5; 11694: data <= 'd5; 11695: data <= 'd1; 11696: data <= 'd1; 11697: data <= 'd1; 11698: data <= 'd1; 11699: data <= 'd1; 11700: data <= 'd5; 11701: data <= 'd5; 11702: data <= 'd2; 11703: data <= 'd0; 11704: data <= 'd0; 11705: data <= 'd0; 11706: data <= 'd0; 11707: data <= 'd0; 11708: data <= 'd0; 11709: data <= 'd0; 11710: data <= 'd0; 11711: data <= 'd0; 11712: data <= 'd0; 11713: data <= 'd0; 11714: data <= 'd0; 11715: data <= 'd0; 11716: data <= 'd0; 11717: data <= 'd0; 11718: data <= 'd0; 11719: data <= 'd0; 11720: data <= 'd2; 11721: data <= 'd1; 11722: data <= 'd5; 11723: data <= 'd5; 11724: data <= 'd3; 11725: data <= 'd6; 11726: data <= 'd6; 11727: data <= 'd6; 11728: data <= 'd6; 11729: data <= 'd6; 11730: data <= 'd6; 11731: data <= 'd6; 11732: data <= 'd6; 11733: data <= 'd3; 11734: data <= 'd5; 11735: data <= 'd2; 11736: data <= 'd0; 11737: data <= 'd0; 11738: data <= 'd0; 11739: data <= 'd0; 11740: data <= 'd0; 11741: data <= 'd0; 11742: data <= 'd0; 11743: data <= 'd0; 11744: data <= 'd0; 11745: data <= 'd0; 11746: data <= 'd0; 11747: data <= 'd0; 11748: data <= 'd0; 11749: data <= 'd0; 11750: data <= 'd0; 11751: data <= 'd0; 11752: data <= 'd2; 11753: data <= 'd5; 11754: data <= 'd3; 11755: data <= 'd6; 11756: data <= 'd3; 11757: data <= 'd1; 11758: data <= 'd1; 11759: data <= 'd1; 11760: data <= 'd1; 11761: data <= 'd1; 11762: data <= 'd1; 11763: data <= 'd1; 11764: data <= 'd1; 11765: data <= 'd1; 11766: data <= 'd3; 11767: data <= 'd2; 11768: data <= 'd0; 11769: data <= 'd0; 11770: data <= 'd0; 11771: data <= 'd0; 11772: data <= 'd0; 11773: data <= 'd0; 11774: data <= 'd0; 11775: data <= 'd0; 11776: data <= 'd0; 11777: data <= 'd0; 11778: data <= 'd0; 11779: data <= 'd0; 11780: data <= 'd0; 11781: data <= 'd0; 11782: data <= 'd0; 11783: data <= 'd0; 11784: data <= 'd2; 11785: data <= 'd5; 11786: data <= 'd3; 11787: data <= 'd1; 11788: data <= 'd1; 11789: data <= 'd1; 11790: data <= 'd5; 11791: data <= 'd5; 11792: data <= 'd5; 11793: data <= 'd5; 11794: data <= 'd5; 11795: data <= 'd5; 11796: data <= 'd5; 11797: data <= 'd1; 11798: data <= 'd1; 11799: data <= 'd2; 11800: data <= 'd0; 11801: data <= 'd0; 11802: data <= 'd0; 11803: data <= 'd0; 11804: data <= 'd0; 11805: data <= 'd0; 11806: data <= 'd0; 11807: data <= 'd0; 11808: data <= 'd0; 11809: data <= 'd0; 11810: data <= 'd0; 11811: data <= 'd0; 11812: data <= 'd0; 11813: data <= 'd0; 11814: data <= 'd0; 11815: data <= 'd0; 11816: data <= 'd2; 11817: data <= 'd6; 11818: data <= 'd1; 11819: data <= 'd5; 11820: data <= 'd2; 11821: data <= 'd2; 11822: data <= 'd2; 11823: data <= 'd2; 11824: data <= 'd2; 11825: data <= 'd2; 11826: data <= 'd2; 11827: data <= 'd2; 11828: data <= 'd2; 11829: data <= 'd2; 11830: data <= 'd5; 11831: data <= 'd2; 11832: data <= 'd0; 11833: data <= 'd0; 11834: data <= 'd0; 11835: data <= 'd0; 11836: data <= 'd0; 11837: data <= 'd0; 11838: data <= 'd0; 11839: data <= 'd0; 11840: data <= 'd0; 11841: data <= 'd0; 11842: data <= 'd0; 11843: data <= 'd0; 11844: data <= 'd0; 11845: data <= 'd0; 11846: data <= 'd2; 11847: data <= 'd2; 11848: data <= 'd2; 11849: data <= 'd1; 11850: data <= 'd5; 11851: data <= 'd2; 11852: data <= 'd8; 11853: data <= 'd8; 11854: data <= 'd8; 11855: data <= 'd8; 11856: data <= 'd8; 11857: data <= 'd9; 11858: data <= 'd9; 11859: data <= 'd8; 11860: data <= 'd8; 11861: data <= 'd8; 11862: data <= 'd2; 11863: data <= 'd2; 11864: data <= 'd0; 11865: data <= 'd0; 11866: data <= 'd0; 11867: data <= 'd0; 11868: data <= 'd0; 11869: data <= 'd0; 11870: data <= 'd0; 11871: data <= 'd0; 11872: data <= 'd0; 11873: data <= 'd0; 11874: data <= 'd0; 11875: data <= 'd0; 11876: data <= 'd0; 11877: data <= 'd0; 11878: data <= 'd2; 11879: data <= 'd1; 11880: data <= 'd2; 11881: data <= 'd1; 11882: data <= 'd2; 11883: data <= 'd8; 11884: data <= 'd8; 11885: data <= 'd9; 11886: data <= 'd9; 11887: data <= 'd2; 11888: data <= 'd9; 11889: data <= 'd11; 11890: data <= 'd11; 11891: data <= 'd10; 11892: data <= 'd2; 11893: data <= 'd9; 11894: data <= 'd2; 11895: data <= 'd2; 11896: data <= 'd0; 11897: data <= 'd0; 11898: data <= 'd0; 11899: data <= 'd0; 11900: data <= 'd0; 11901: data <= 'd0; 11902: data <= 'd0; 11903: data <= 'd0; 11904: data <= 'd0; 11905: data <= 'd0; 11906: data <= 'd0; 11907: data <= 'd0; 11908: data <= 'd0; 11909: data <= 'd0; 11910: data <= 'd2; 11911: data <= 'd5; 11912: data <= 'd1; 11913: data <= 'd2; 11914: data <= 'd9; 11915: data <= 'd10; 11916: data <= 'd9; 11917: data <= 'd9; 11918: data <= 'd10; 11919: data <= 'd11; 11920: data <= 'd10; 11921: data <= 'd11; 11922: data <= 'd11; 11923: data <= 'd10; 11924: data <= 'd11; 11925: data <= 'd10; 11926: data <= 'd9; 11927: data <= 'd2; 11928: data <= 'd0; 11929: data <= 'd0; 11930: data <= 'd0; 11931: data <= 'd0; 11932: data <= 'd0; 11933: data <= 'd0; 11934: data <= 'd0; 11935: data <= 'd0; 11936: data <= 'd0; 11937: data <= 'd0; 11938: data <= 'd0; 11939: data <= 'd0; 11940: data <= 'd0; 11941: data <= 'd0; 11942: data <= 'd0; 11943: data <= 'd2; 11944: data <= 'd5; 11945: data <= 'd5; 11946: data <= 'd2; 11947: data <= 'd8; 11948: data <= 'd9; 11949: data <= 'd9; 11950: data <= 'd10; 11951: data <= 'd10; 11952: data <= 'd10; 11953: data <= 'd8; 11954: data <= 'd8; 11955: data <= 'd10; 11956: data <= 'd10; 11957: data <= 'd9; 11958: data <= 'd2; 11959: data <= 'd0; 11960: data <= 'd0; 11961: data <= 'd0; 11962: data <= 'd0; 11963: data <= 'd0; 11964: data <= 'd0; 11965: data <= 'd0; 11966: data <= 'd0; 11967: data <= 'd0; 11968: data <= 'd0; 11969: data <= 'd0; 11970: data <= 'd0; 11971: data <= 'd0; 11972: data <= 'd0; 11973: data <= 'd0; 11974: data <= 'd0; 11975: data <= 'd0; 11976: data <= 'd2; 11977: data <= 'd2; 11978: data <= 'd2; 11979: data <= 'd8; 11980: data <= 'd8; 11981: data <= 'd9; 11982: data <= 'd9; 11983: data <= 'd10; 11984: data <= 'd10; 11985: data <= 'd9; 11986: data <= 'd9; 11987: data <= 'd10; 11988: data <= 'd10; 11989: data <= 'd9; 11990: data <= 'd2; 11991: data <= 'd0; 11992: data <= 'd0; 11993: data <= 'd0; 11994: data <= 'd0; 11995: data <= 'd0; 11996: data <= 'd0; 11997: data <= 'd0; 11998: data <= 'd0; 11999: data <= 'd0; 12000: data <= 'd0; 12001: data <= 'd0; 12002: data <= 'd0; 12003: data <= 'd0; 12004: data <= 'd0; 12005: data <= 'd0; 12006: data <= 'd0; 12007: data <= 'd0; 12008: data <= 'd0; 12009: data <= 'd0; 12010: data <= 'd0; 12011: data <= 'd2; 12012: data <= 'd5; 12013: data <= 'd5; 12014: data <= 'd8; 12015: data <= 'd9; 12016: data <= 'd9; 12017: data <= 'd9; 12018: data <= 'd9; 12019: data <= 'd9; 12020: data <= 'd9; 12021: data <= 'd5; 12022: data <= 'd2; 12023: data <= 'd0; 12024: data <= 'd0; 12025: data <= 'd0; 12026: data <= 'd0; 12027: data <= 'd0; 12028: data <= 'd0; 12029: data <= 'd0; 12030: data <= 'd0; 12031: data <= 'd0; 12032: data <= 'd0; 12033: data <= 'd0; 12034: data <= 'd0; 12035: data <= 'd0; 12036: data <= 'd0; 12037: data <= 'd0; 12038: data <= 'd0; 12039: data <= 'd0; 12040: data <= 'd0; 12041: data <= 'd0; 12042: data <= 'd2; 12043: data <= 'd1; 12044: data <= 'd1; 12045: data <= 'd1; 12046: data <= 'd3; 12047: data <= 'd3; 12048: data <= 'd3; 12049: data <= 'd5; 12050: data <= 'd5; 12051: data <= 'd3; 12052: data <= 'd3; 12053: data <= 'd1; 12054: data <= 'd2; 12055: data <= 'd0; 12056: data <= 'd0; 12057: data <= 'd0; 12058: data <= 'd0; 12059: data <= 'd0; 12060: data <= 'd0; 12061: data <= 'd0; 12062: data <= 'd0; 12063: data <= 'd0; 12064: data <= 'd0; 12065: data <= 'd0; 12066: data <= 'd0; 12067: data <= 'd0; 12068: data <= 'd0; 12069: data <= 'd0; 12070: data <= 'd0; 12071: data <= 'd0; 12072: data <= 'd0; 12073: data <= 'd0; 12074: data <= 'd2; 12075: data <= 'd7; 12076: data <= 'd1; 12077: data <= 'd5; 12078: data <= 'd2; 12079: data <= 'd3; 12080: data <= 'd3; 12081: data <= 'd1; 12082: data <= 'd1; 12083: data <= 'd3; 12084: data <= 'd3; 12085: data <= 'd1; 12086: data <= 'd2; 12087: data <= 'd0; 12088: data <= 'd0; 12089: data <= 'd0; 12090: data <= 'd0; 12091: data <= 'd0; 12092: data <= 'd0; 12093: data <= 'd0; 12094: data <= 'd0; 12095: data <= 'd0; 12096: data <= 'd0; 12097: data <= 'd0; 12098: data <= 'd0; 12099: data <= 'd0; 12100: data <= 'd0; 12101: data <= 'd0; 12102: data <= 'd0; 12103: data <= 'd0; 12104: data <= 'd0; 12105: data <= 'd0; 12106: data <= 'd2; 12107: data <= 'd8; 12108: data <= 'd9; 12109: data <= 'd10; 12110: data <= 'd10; 12111: data <= 'd2; 12112: data <= 'd3; 12113: data <= 'd1; 12114: data <= 'd1; 12115: data <= 'd3; 12116: data <= 'd1; 12117: data <= 'd1; 12118: data <= 'd2; 12119: data <= 'd0; 12120: data <= 'd0; 12121: data <= 'd0; 12122: data <= 'd0; 12123: data <= 'd0; 12124: data <= 'd0; 12125: data <= 'd0; 12126: data <= 'd0; 12127: data <= 'd0; 12128: data <= 'd0; 12129: data <= 'd0; 12130: data <= 'd0; 12131: data <= 'd0; 12132: data <= 'd0; 12133: data <= 'd0; 12134: data <= 'd0; 12135: data <= 'd0; 12136: data <= 'd0; 12137: data <= 'd0; 12138: data <= 'd0; 12139: data <= 'd2; 12140: data <= 'd8; 12141: data <= 'd9; 12142: data <= 'd9; 12143: data <= 'd2; 12144: data <= 'd5; 12145: data <= 'd5; 12146: data <= 'd5; 12147: data <= 'd2; 12148: data <= 'd2; 12149: data <= 'd2; 12150: data <= 'd2; 12151: data <= 'd0; 12152: data <= 'd0; 12153: data <= 'd0; 12154: data <= 'd0; 12155: data <= 'd0; 12156: data <= 'd0; 12157: data <= 'd0; 12158: data <= 'd0; 12159: data <= 'd0; 12160: data <= 'd0; 12161: data <= 'd0; 12162: data <= 'd0; 12163: data <= 'd0; 12164: data <= 'd0; 12165: data <= 'd0; 12166: data <= 'd0; 12167: data <= 'd0; 12168: data <= 'd0; 12169: data <= 'd0; 12170: data <= 'd0; 12171: data <= 'd2; 12172: data <= 'd2; 12173: data <= 'd2; 12174: data <= 'd2; 12175: data <= 'd3; 12176: data <= 'd3; 12177: data <= 'd1; 12178: data <= 'd3; 12179: data <= 'd3; 12180: data <= 'd3; 12181: data <= 'd5; 12182: data <= 'd0; 12183: data <= 'd0; 12184: data <= 'd0; 12185: data <= 'd0; 12186: data <= 'd0; 12187: data <= 'd0; 12188: data <= 'd0; 12189: data <= 'd0; 12190: data <= 'd0; 12191: data <= 'd0; 12192: data <= 'd0; 12193: data <= 'd0; 12194: data <= 'd0; 12195: data <= 'd0; 12196: data <= 'd0; 12197: data <= 'd0; 12198: data <= 'd0; 12199: data <= 'd0; 12200: data <= 'd0; 12201: data <= 'd0; 12202: data <= 'd0; 12203: data <= 'd2; 12204: data <= 'd4; 12205: data <= 'd7; 12206: data <= 'd7; 12207: data <= 'd2; 12208: data <= 'd2; 12209: data <= 'd2; 12210: data <= 'd5; 12211: data <= 'd5; 12212: data <= 'd4; 12213: data <= 'd2; 12214: data <= 'd0; 12215: data <= 'd0; 12216: data <= 'd0; 12217: data <= 'd0; 12218: data <= 'd0; 12219: data <= 'd0; 12220: data <= 'd0; 12221: data <= 'd0; 12222: data <= 'd0; 12223: data <= 'd0; 12224: data <= 'd0; 12225: data <= 'd0; 12226: data <= 'd0; 12227: data <= 'd0; 12228: data <= 'd0; 12229: data <= 'd0; 12230: data <= 'd0; 12231: data <= 'd0; 12232: data <= 'd0; 12233: data <= 'd0; 12234: data <= 'd0; 12235: data <= 'd2; 12236: data <= 'd4; 12237: data <= 'd7; 12238: data <= 'd2; 12239: data <= 'd0; 12240: data <= 'd0; 12241: data <= 'd0; 12242: data <= 'd2; 12243: data <= 'd4; 12244: data <= 'd4; 12245: data <= 'd2; 12246: data <= 'd0; 12247: data <= 'd0; 12248: data <= 'd0; 12249: data <= 'd0; 12250: data <= 'd0; 12251: data <= 'd0; 12252: data <= 'd0; 12253: data <= 'd0; 12254: data <= 'd0; 12255: data <= 'd0; 12256: data <= 'd0; 12257: data <= 'd0; 12258: data <= 'd0; 12259: data <= 'd0; 12260: data <= 'd0; 12261: data <= 'd0; 12262: data <= 'd0; 12263: data <= 'd0; 12264: data <= 'd0; 12265: data <= 'd0; 12266: data <= 'd0; 12267: data <= 'd2; 12268: data <= 'd2; 12269: data <= 'd2; 12270: data <= 'd0; 12271: data <= 'd0; 12272: data <= 'd0; 12273: data <= 'd0; 12274: data <= 'd2; 12275: data <= 'd2; 12276: data <= 'd2; 12277: data <= 'd0; 12278: data <= 'd0; 12279: data <= 'd0; 12280: data <= 'd0; 12281: data <= 'd0; 12282: data <= 'd0; 12283: data <= 'd0; 12284: data <= 'd0; 12285: data <= 'd0; 12286: data <= 'd0; 12287: data <= 'd0; 12288: data <= 'd0; 12289: data <= 'd0; 12290: data <= 'd0; 12291: data <= 'd0; 12292: data <= 'd0; 12293: data <= 'd0; 12294: data <= 'd0; 12295: data <= 'd0; 12296: data <= 'd0; 12297: data <= 'd0; 12298: data <= 'd0; 12299: data <= 'd0; 12300: data <= 'd0; 12301: data <= 'd0; 12302: data <= 'd0; 12303: data <= 'd0; 12304: data <= 'd0; 12305: data <= 'd0; 12306: data <= 'd0; 12307: data <= 'd0; 12308: data <= 'd0; 12309: data <= 'd0; 12310: data <= 'd0; 12311: data <= 'd0; 12312: data <= 'd0; 12313: data <= 'd0; 12314: data <= 'd0; 12315: data <= 'd0; 12316: data <= 'd0; 12317: data <= 'd0; 12318: data <= 'd0; 12319: data <= 'd0; 12320: data <= 'd0; 12321: data <= 'd0; 12322: data <= 'd0; 12323: data <= 'd0; 12324: data <= 'd0; 12325: data <= 'd0; 12326: data <= 'd0; 12327: data <= 'd0; 12328: data <= 'd0; 12329: data <= 'd0; 12330: data <= 'd0; 12331: data <= 'd0; 12332: data <= 'd0; 12333: data <= 'd0; 12334: data <= 'd0; 12335: data <= 'd0; 12336: data <= 'd0; 12337: data <= 'd0; 12338: data <= 'd0; 12339: data <= 'd0; 12340: data <= 'd0; 12341: data <= 'd0; 12342: data <= 'd0; 12343: data <= 'd0; 12344: data <= 'd0; 12345: data <= 'd0; 12346: data <= 'd0; 12347: data <= 'd0; 12348: data <= 'd0; 12349: data <= 'd0; 12350: data <= 'd0; 12351: data <= 'd0; 12352: data <= 'd0; 12353: data <= 'd0; 12354: data <= 'd0; 12355: data <= 'd0; 12356: data <= 'd0; 12357: data <= 'd0; 12358: data <= 'd0; 12359: data <= 'd0; 12360: data <= 'd0; 12361: data <= 'd0; 12362: data <= 'd0; 12363: data <= 'd0; 12364: data <= 'd0; 12365: data <= 'd0; 12366: data <= 'd0; 12367: data <= 'd0; 12368: data <= 'd0; 12369: data <= 'd0; 12370: data <= 'd0; 12371: data <= 'd0; 12372: data <= 'd0; 12373: data <= 'd0; 12374: data <= 'd0; 12375: data <= 'd0; 12376: data <= 'd0; 12377: data <= 'd0; 12378: data <= 'd0; 12379: data <= 'd0; 12380: data <= 'd0; 12381: data <= 'd0; 12382: data <= 'd0; 12383: data <= 'd0; 12384: data <= 'd0; 12385: data <= 'd0; 12386: data <= 'd0; 12387: data <= 'd0; 12388: data <= 'd0; 12389: data <= 'd0; 12390: data <= 'd0; 12391: data <= 'd0; 12392: data <= 'd0; 12393: data <= 'd0; 12394: data <= 'd0; 12395: data <= 'd0; 12396: data <= 'd0; 12397: data <= 'd0; 12398: data <= 'd0; 12399: data <= 'd0; 12400: data <= 'd0; 12401: data <= 'd0; 12402: data <= 'd0; 12403: data <= 'd0; 12404: data <= 'd0; 12405: data <= 'd0; 12406: data <= 'd0; 12407: data <= 'd0; 12408: data <= 'd0; 12409: data <= 'd0; 12410: data <= 'd0; 12411: data <= 'd0; 12412: data <= 'd0; 12413: data <= 'd0; 12414: data <= 'd0; 12415: data <= 'd0; 12416: data <= 'd0; 12417: data <= 'd0; 12418: data <= 'd0; 12419: data <= 'd0; 12420: data <= 'd0; 12421: data <= 'd0; 12422: data <= 'd0; 12423: data <= 'd0; 12424: data <= 'd0; 12425: data <= 'd0; 12426: data <= 'd0; 12427: data <= 'd0; 12428: data <= 'd0; 12429: data <= 'd0; 12430: data <= 'd0; 12431: data <= 'd0; 12432: data <= 'd0; 12433: data <= 'd0; 12434: data <= 'd0; 12435: data <= 'd0; 12436: data <= 'd0; 12437: data <= 'd0; 12438: data <= 'd0; 12439: data <= 'd0; 12440: data <= 'd0; 12441: data <= 'd0; 12442: data <= 'd0; 12443: data <= 'd0; 12444: data <= 'd0; 12445: data <= 'd0; 12446: data <= 'd0; 12447: data <= 'd0; 12448: data <= 'd0; 12449: data <= 'd0; 12450: data <= 'd0; 12451: data <= 'd0; 12452: data <= 'd0; 12453: data <= 'd0; 12454: data <= 'd0; 12455: data <= 'd0; 12456: data <= 'd0; 12457: data <= 'd0; 12458: data <= 'd0; 12459: data <= 'd0; 12460: data <= 'd0; 12461: data <= 'd0; 12462: data <= 'd0; 12463: data <= 'd0; 12464: data <= 'd0; 12465: data <= 'd0; 12466: data <= 'd0; 12467: data <= 'd0; 12468: data <= 'd0; 12469: data <= 'd0; 12470: data <= 'd0; 12471: data <= 'd0; 12472: data <= 'd0; 12473: data <= 'd0; 12474: data <= 'd0; 12475: data <= 'd0; 12476: data <= 'd0; 12477: data <= 'd0; 12478: data <= 'd0; 12479: data <= 'd0; 12480: data <= 'd0; 12481: data <= 'd0; 12482: data <= 'd0; 12483: data <= 'd0; 12484: data <= 'd0; 12485: data <= 'd0; 12486: data <= 'd0; 12487: data <= 'd0; 12488: data <= 'd0; 12489: data <= 'd0; 12490: data <= 'd0; 12491: data <= 'd0; 12492: data <= 'd0; 12493: data <= 'd0; 12494: data <= 'd0; 12495: data <= 'd0; 12496: data <= 'd0; 12497: data <= 'd0; 12498: data <= 'd0; 12499: data <= 'd0; 12500: data <= 'd0; 12501: data <= 'd0; 12502: data <= 'd0; 12503: data <= 'd0; 12504: data <= 'd0; 12505: data <= 'd0; 12506: data <= 'd0; 12507: data <= 'd0; 12508: data <= 'd0; 12509: data <= 'd0; 12510: data <= 'd0; 12511: data <= 'd0; 12512: data <= 'd0; 12513: data <= 'd0; 12514: data <= 'd0; 12515: data <= 'd0; 12516: data <= 'd0; 12517: data <= 'd0; 12518: data <= 'd0; 12519: data <= 'd0; 12520: data <= 'd0; 12521: data <= 'd0; 12522: data <= 'd0; 12523: data <= 'd0; 12524: data <= 'd0; 12525: data <= 'd0; 12526: data <= 'd0; 12527: data <= 'd0; 12528: data <= 'd0; 12529: data <= 'd0; 12530: data <= 'd0; 12531: data <= 'd0; 12532: data <= 'd0; 12533: data <= 'd0; 12534: data <= 'd0; 12535: data <= 'd0; 12536: data <= 'd0; 12537: data <= 'd0; 12538: data <= 'd0; 12539: data <= 'd0; 12540: data <= 'd0; 12541: data <= 'd0; 12542: data <= 'd0; 12543: data <= 'd0; 12544: data <= 'd0; 12545: data <= 'd0; 12546: data <= 'd0; 12547: data <= 'd0; 12548: data <= 'd0; 12549: data <= 'd0; 12550: data <= 'd0; 12551: data <= 'd0; 12552: data <= 'd0; 12553: data <= 'd0; 12554: data <= 'd0; 12555: data <= 'd0; 12556: data <= 'd0; 12557: data <= 'd0; 12558: data <= 'd0; 12559: data <= 'd0; 12560: data <= 'd0; 12561: data <= 'd0; 12562: data <= 'd0; 12563: data <= 'd0; 12564: data <= 'd0; 12565: data <= 'd0; 12566: data <= 'd0; 12567: data <= 'd0; 12568: data <= 'd0; 12569: data <= 'd0; 12570: data <= 'd0; 12571: data <= 'd0; 12572: data <= 'd0; 12573: data <= 'd0; 12574: data <= 'd0; 12575: data <= 'd0; 12576: data <= 'd0; 12577: data <= 'd0; 12578: data <= 'd0; 12579: data <= 'd0; 12580: data <= 'd0; 12581: data <= 'd0; 12582: data <= 'd0; 12583: data <= 'd0; 12584: data <= 'd0; 12585: data <= 'd0; 12586: data <= 'd0; 12587: data <= 'd0; 12588: data <= 'd0; 12589: data <= 'd2; 12590: data <= 'd2; 12591: data <= 'd2; 12592: data <= 'd2; 12593: data <= 'd2; 12594: data <= 'd2; 12595: data <= 'd0; 12596: data <= 'd0; 12597: data <= 'd0; 12598: data <= 'd0; 12599: data <= 'd0; 12600: data <= 'd0; 12601: data <= 'd0; 12602: data <= 'd0; 12603: data <= 'd0; 12604: data <= 'd0; 12605: data <= 'd0; 12606: data <= 'd0; 12607: data <= 'd0; 12608: data <= 'd0; 12609: data <= 'd0; 12610: data <= 'd0; 12611: data <= 'd0; 12612: data <= 'd0; 12613: data <= 'd0; 12614: data <= 'd0; 12615: data <= 'd0; 12616: data <= 'd0; 12617: data <= 'd0; 12618: data <= 'd0; 12619: data <= 'd2; 12620: data <= 'd2; 12621: data <= 'd6; 12622: data <= 'd6; 12623: data <= 'd6; 12624: data <= 'd6; 12625: data <= 'd6; 12626: data <= 'd6; 12627: data <= 'd2; 12628: data <= 'd2; 12629: data <= 'd0; 12630: data <= 'd0; 12631: data <= 'd0; 12632: data <= 'd0; 12633: data <= 'd0; 12634: data <= 'd0; 12635: data <= 'd0; 12636: data <= 'd0; 12637: data <= 'd0; 12638: data <= 'd0; 12639: data <= 'd0; 12640: data <= 'd0; 12641: data <= 'd0; 12642: data <= 'd0; 12643: data <= 'd0; 12644: data <= 'd0; 12645: data <= 'd0; 12646: data <= 'd0; 12647: data <= 'd0; 12648: data <= 'd0; 12649: data <= 'd0; 12650: data <= 'd2; 12651: data <= 'd1; 12652: data <= 'd3; 12653: data <= 'd6; 12654: data <= 'd6; 12655: data <= 'd6; 12656: data <= 'd6; 12657: data <= 'd6; 12658: data <= 'd6; 12659: data <= 'd6; 12660: data <= 'd3; 12661: data <= 'd2; 12662: data <= 'd0; 12663: data <= 'd0; 12664: data <= 'd0; 12665: data <= 'd0; 12666: data <= 'd0; 12667: data <= 'd0; 12668: data <= 'd0; 12669: data <= 'd0; 12670: data <= 'd0; 12671: data <= 'd0; 12672: data <= 'd0; 12673: data <= 'd0; 12674: data <= 'd0; 12675: data <= 'd0; 12676: data <= 'd0; 12677: data <= 'd0; 12678: data <= 'd0; 12679: data <= 'd0; 12680: data <= 'd0; 12681: data <= 'd2; 12682: data <= 'd1; 12683: data <= 'd1; 12684: data <= 'd1; 12685: data <= 'd3; 12686: data <= 'd6; 12687: data <= 'd6; 12688: data <= 'd6; 12689: data <= 'd6; 12690: data <= 'd6; 12691: data <= 'd3; 12692: data <= 'd1; 12693: data <= 'd1; 12694: data <= 'd2; 12695: data <= 'd0; 12696: data <= 'd0; 12697: data <= 'd0; 12698: data <= 'd0; 12699: data <= 'd0; 12700: data <= 'd0; 12701: data <= 'd0; 12702: data <= 'd0; 12703: data <= 'd0; 12704: data <= 'd0; 12705: data <= 'd0; 12706: data <= 'd0; 12707: data <= 'd0; 12708: data <= 'd0; 12709: data <= 'd0; 12710: data <= 'd0; 12711: data <= 'd0; 12712: data <= 'd0; 12713: data <= 'd2; 12714: data <= 'd1; 12715: data <= 'd1; 12716: data <= 'd5; 12717: data <= 'd5; 12718: data <= 'd5; 12719: data <= 'd1; 12720: data <= 'd1; 12721: data <= 'd1; 12722: data <= 'd1; 12723: data <= 'd1; 12724: data <= 'd5; 12725: data <= 'd5; 12726: data <= 'd2; 12727: data <= 'd0; 12728: data <= 'd0; 12729: data <= 'd0; 12730: data <= 'd0; 12731: data <= 'd0; 12732: data <= 'd0; 12733: data <= 'd0; 12734: data <= 'd0; 12735: data <= 'd0; 12736: data <= 'd0; 12737: data <= 'd0; 12738: data <= 'd0; 12739: data <= 'd0; 12740: data <= 'd0; 12741: data <= 'd0; 12742: data <= 'd0; 12743: data <= 'd0; 12744: data <= 'd2; 12745: data <= 'd1; 12746: data <= 'd5; 12747: data <= 'd5; 12748: data <= 'd3; 12749: data <= 'd6; 12750: data <= 'd6; 12751: data <= 'd6; 12752: data <= 'd6; 12753: data <= 'd6; 12754: data <= 'd6; 12755: data <= 'd6; 12756: data <= 'd6; 12757: data <= 'd3; 12758: data <= 'd5; 12759: data <= 'd2; 12760: data <= 'd0; 12761: data <= 'd0; 12762: data <= 'd0; 12763: data <= 'd0; 12764: data <= 'd0; 12765: data <= 'd0; 12766: data <= 'd0; 12767: data <= 'd0; 12768: data <= 'd0; 12769: data <= 'd0; 12770: data <= 'd0; 12771: data <= 'd0; 12772: data <= 'd0; 12773: data <= 'd0; 12774: data <= 'd0; 12775: data <= 'd0; 12776: data <= 'd2; 12777: data <= 'd5; 12778: data <= 'd3; 12779: data <= 'd6; 12780: data <= 'd3; 12781: data <= 'd1; 12782: data <= 'd1; 12783: data <= 'd1; 12784: data <= 'd1; 12785: data <= 'd1; 12786: data <= 'd1; 12787: data <= 'd1; 12788: data <= 'd1; 12789: data <= 'd1; 12790: data <= 'd3; 12791: data <= 'd2; 12792: data <= 'd0; 12793: data <= 'd0; 12794: data <= 'd0; 12795: data <= 'd0; 12796: data <= 'd0; 12797: data <= 'd0; 12798: data <= 'd0; 12799: data <= 'd0; 12800: data <= 'd0; 12801: data <= 'd0; 12802: data <= 'd0; 12803: data <= 'd0; 12804: data <= 'd0; 12805: data <= 'd0; 12806: data <= 'd0; 12807: data <= 'd0; 12808: data <= 'd2; 12809: data <= 'd5; 12810: data <= 'd3; 12811: data <= 'd1; 12812: data <= 'd1; 12813: data <= 'd1; 12814: data <= 'd5; 12815: data <= 'd5; 12816: data <= 'd5; 12817: data <= 'd5; 12818: data <= 'd5; 12819: data <= 'd5; 12820: data <= 'd5; 12821: data <= 'd1; 12822: data <= 'd1; 12823: data <= 'd2; 12824: data <= 'd0; 12825: data <= 'd0; 12826: data <= 'd0; 12827: data <= 'd0; 12828: data <= 'd0; 12829: data <= 'd0; 12830: data <= 'd0; 12831: data <= 'd0; 12832: data <= 'd0; 12833: data <= 'd0; 12834: data <= 'd0; 12835: data <= 'd0; 12836: data <= 'd0; 12837: data <= 'd0; 12838: data <= 'd0; 12839: data <= 'd0; 12840: data <= 'd2; 12841: data <= 'd6; 12842: data <= 'd1; 12843: data <= 'd5; 12844: data <= 'd2; 12845: data <= 'd2; 12846: data <= 'd2; 12847: data <= 'd2; 12848: data <= 'd2; 12849: data <= 'd2; 12850: data <= 'd2; 12851: data <= 'd2; 12852: data <= 'd2; 12853: data <= 'd2; 12854: data <= 'd5; 12855: data <= 'd2; 12856: data <= 'd0; 12857: data <= 'd0; 12858: data <= 'd0; 12859: data <= 'd0; 12860: data <= 'd0; 12861: data <= 'd0; 12862: data <= 'd0; 12863: data <= 'd0; 12864: data <= 'd0; 12865: data <= 'd0; 12866: data <= 'd0; 12867: data <= 'd0; 12868: data <= 'd0; 12869: data <= 'd0; 12870: data <= 'd2; 12871: data <= 'd2; 12872: data <= 'd2; 12873: data <= 'd1; 12874: data <= 'd5; 12875: data <= 'd2; 12876: data <= 'd8; 12877: data <= 'd8; 12878: data <= 'd8; 12879: data <= 'd8; 12880: data <= 'd8; 12881: data <= 'd9; 12882: data <= 'd9; 12883: data <= 'd8; 12884: data <= 'd8; 12885: data <= 'd8; 12886: data <= 'd2; 12887: data <= 'd2; 12888: data <= 'd0; 12889: data <= 'd0; 12890: data <= 'd0; 12891: data <= 'd0; 12892: data <= 'd0; 12893: data <= 'd0; 12894: data <= 'd0; 12895: data <= 'd0; 12896: data <= 'd0; 12897: data <= 'd0; 12898: data <= 'd0; 12899: data <= 'd0; 12900: data <= 'd0; 12901: data <= 'd0; 12902: data <= 'd2; 12903: data <= 'd1; 12904: data <= 'd2; 12905: data <= 'd1; 12906: data <= 'd2; 12907: data <= 'd8; 12908: data <= 'd8; 12909: data <= 'd9; 12910: data <= 'd9; 12911: data <= 'd2; 12912: data <= 'd9; 12913: data <= 'd11; 12914: data <= 'd11; 12915: data <= 'd10; 12916: data <= 'd2; 12917: data <= 'd9; 12918: data <= 'd2; 12919: data <= 'd2; 12920: data <= 'd0; 12921: data <= 'd0; 12922: data <= 'd0; 12923: data <= 'd0; 12924: data <= 'd0; 12925: data <= 'd0; 12926: data <= 'd0; 12927: data <= 'd0; 12928: data <= 'd0; 12929: data <= 'd0; 12930: data <= 'd0; 12931: data <= 'd0; 12932: data <= 'd0; 12933: data <= 'd0; 12934: data <= 'd2; 12935: data <= 'd5; 12936: data <= 'd1; 12937: data <= 'd2; 12938: data <= 'd9; 12939: data <= 'd10; 12940: data <= 'd9; 12941: data <= 'd9; 12942: data <= 'd10; 12943: data <= 'd11; 12944: data <= 'd10; 12945: data <= 'd11; 12946: data <= 'd11; 12947: data <= 'd10; 12948: data <= 'd11; 12949: data <= 'd10; 12950: data <= 'd9; 12951: data <= 'd2; 12952: data <= 'd0; 12953: data <= 'd0; 12954: data <= 'd0; 12955: data <= 'd0; 12956: data <= 'd0; 12957: data <= 'd0; 12958: data <= 'd0; 12959: data <= 'd0; 12960: data <= 'd0; 12961: data <= 'd0; 12962: data <= 'd0; 12963: data <= 'd0; 12964: data <= 'd0; 12965: data <= 'd0; 12966: data <= 'd0; 12967: data <= 'd2; 12968: data <= 'd5; 12969: data <= 'd5; 12970: data <= 'd2; 12971: data <= 'd8; 12972: data <= 'd9; 12973: data <= 'd9; 12974: data <= 'd10; 12975: data <= 'd10; 12976: data <= 'd10; 12977: data <= 'd8; 12978: data <= 'd8; 12979: data <= 'd10; 12980: data <= 'd10; 12981: data <= 'd9; 12982: data <= 'd2; 12983: data <= 'd0; 12984: data <= 'd0; 12985: data <= 'd0; 12986: data <= 'd0; 12987: data <= 'd0; 12988: data <= 'd0; 12989: data <= 'd0; 12990: data <= 'd0; 12991: data <= 'd0; 12992: data <= 'd0; 12993: data <= 'd0; 12994: data <= 'd0; 12995: data <= 'd0; 12996: data <= 'd0; 12997: data <= 'd0; 12998: data <= 'd0; 12999: data <= 'd0; 13000: data <= 'd2; 13001: data <= 'd2; 13002: data <= 'd2; 13003: data <= 'd8; 13004: data <= 'd8; 13005: data <= 'd9; 13006: data <= 'd9; 13007: data <= 'd10; 13008: data <= 'd10; 13009: data <= 'd9; 13010: data <= 'd9; 13011: data <= 'd10; 13012: data <= 'd10; 13013: data <= 'd9; 13014: data <= 'd2; 13015: data <= 'd0; 13016: data <= 'd0; 13017: data <= 'd0; 13018: data <= 'd0; 13019: data <= 'd0; 13020: data <= 'd0; 13021: data <= 'd0; 13022: data <= 'd0; 13023: data <= 'd0; 13024: data <= 'd0; 13025: data <= 'd0; 13026: data <= 'd0; 13027: data <= 'd0; 13028: data <= 'd0; 13029: data <= 'd0; 13030: data <= 'd0; 13031: data <= 'd0; 13032: data <= 'd0; 13033: data <= 'd0; 13034: data <= 'd2; 13035: data <= 'd2; 13036: data <= 'd5; 13037: data <= 'd5; 13038: data <= 'd8; 13039: data <= 'd9; 13040: data <= 'd9; 13041: data <= 'd9; 13042: data <= 'd9; 13043: data <= 'd9; 13044: data <= 'd9; 13045: data <= 'd5; 13046: data <= 'd2; 13047: data <= 'd0; 13048: data <= 'd0; 13049: data <= 'd0; 13050: data <= 'd0; 13051: data <= 'd0; 13052: data <= 'd0; 13053: data <= 'd0; 13054: data <= 'd0; 13055: data <= 'd0; 13056: data <= 'd0; 13057: data <= 'd0; 13058: data <= 'd0; 13059: data <= 'd0; 13060: data <= 'd0; 13061: data <= 'd0; 13062: data <= 'd0; 13063: data <= 'd0; 13064: data <= 'd0; 13065: data <= 'd2; 13066: data <= 'd7; 13067: data <= 'd1; 13068: data <= 'd1; 13069: data <= 'd1; 13070: data <= 'd3; 13071: data <= 'd3; 13072: data <= 'd3; 13073: data <= 'd5; 13074: data <= 'd5; 13075: data <= 'd3; 13076: data <= 'd3; 13077: data <= 'd1; 13078: data <= 'd2; 13079: data <= 'd0; 13080: data <= 'd0; 13081: data <= 'd0; 13082: data <= 'd0; 13083: data <= 'd0; 13084: data <= 'd0; 13085: data <= 'd0; 13086: data <= 'd0; 13087: data <= 'd0; 13088: data <= 'd0; 13089: data <= 'd0; 13090: data <= 'd0; 13091: data <= 'd0; 13092: data <= 'd0; 13093: data <= 'd0; 13094: data <= 'd0; 13095: data <= 'd0; 13096: data <= 'd0; 13097: data <= 'd2; 13098: data <= 'd7; 13099: data <= 'd7; 13100: data <= 'd5; 13101: data <= 'd1; 13102: data <= 'd3; 13103: data <= 'd3; 13104: data <= 'd3; 13105: data <= 'd1; 13106: data <= 'd1; 13107: data <= 'd3; 13108: data <= 'd3; 13109: data <= 'd1; 13110: data <= 'd2; 13111: data <= 'd0; 13112: data <= 'd0; 13113: data <= 'd0; 13114: data <= 'd0; 13115: data <= 'd0; 13116: data <= 'd0; 13117: data <= 'd0; 13118: data <= 'd0; 13119: data <= 'd0; 13120: data <= 'd0; 13121: data <= 'd0; 13122: data <= 'd0; 13123: data <= 'd0; 13124: data <= 'd0; 13125: data <= 'd0; 13126: data <= 'd0; 13127: data <= 'd0; 13128: data <= 'd0; 13129: data <= 'd0; 13130: data <= 'd2; 13131: data <= 'd9; 13132: data <= 'd9; 13133: data <= 'd2; 13134: data <= 'd1; 13135: data <= 'd3; 13136: data <= 'd3; 13137: data <= 'd1; 13138: data <= 'd1; 13139: data <= 'd3; 13140: data <= 'd1; 13141: data <= 'd1; 13142: data <= 'd8; 13143: data <= 'd2; 13144: data <= 'd0; 13145: data <= 'd0; 13146: data <= 'd0; 13147: data <= 'd0; 13148: data <= 'd0; 13149: data <= 'd0; 13150: data <= 'd0; 13151: data <= 'd0; 13152: data <= 'd0; 13153: data <= 'd0; 13154: data <= 'd0; 13155: data <= 'd0; 13156: data <= 'd0; 13157: data <= 'd0; 13158: data <= 'd0; 13159: data <= 'd0; 13160: data <= 'd0; 13161: data <= 'd0; 13162: data <= 'd2; 13163: data <= 'd9; 13164: data <= 'd9; 13165: data <= 'd2; 13166: data <= 'd2; 13167: data <= 'd2; 13168: data <= 'd5; 13169: data <= 'd5; 13170: data <= 'd5; 13171: data <= 'd2; 13172: data <= 'd2; 13173: data <= 'd2; 13174: data <= 'd8; 13175: data <= 'd2; 13176: data <= 'd0; 13177: data <= 'd0; 13178: data <= 'd0; 13179: data <= 'd0; 13180: data <= 'd0; 13181: data <= 'd0; 13182: data <= 'd0; 13183: data <= 'd0; 13184: data <= 'd0; 13185: data <= 'd0; 13186: data <= 'd0; 13187: data <= 'd0; 13188: data <= 'd0; 13189: data <= 'd0; 13190: data <= 'd0; 13191: data <= 'd0; 13192: data <= 'd0; 13193: data <= 'd0; 13194: data <= 'd0; 13195: data <= 'd2; 13196: data <= 'd2; 13197: data <= 'd1; 13198: data <= 'd3; 13199: data <= 'd3; 13200: data <= 'd3; 13201: data <= 'd1; 13202: data <= 'd3; 13203: data <= 'd3; 13204: data <= 'd3; 13205: data <= 'd5; 13206: data <= 'd2; 13207: data <= 'd0; 13208: data <= 'd0; 13209: data <= 'd0; 13210: data <= 'd0; 13211: data <= 'd0; 13212: data <= 'd0; 13213: data <= 'd0; 13214: data <= 'd0; 13215: data <= 'd0; 13216: data <= 'd0; 13217: data <= 'd0; 13218: data <= 'd0; 13219: data <= 'd0; 13220: data <= 'd0; 13221: data <= 'd0; 13222: data <= 'd0; 13223: data <= 'd0; 13224: data <= 'd0; 13225: data <= 'd0; 13226: data <= 'd0; 13227: data <= 'd2; 13228: data <= 'd4; 13229: data <= 'd7; 13230: data <= 'd7; 13231: data <= 'd2; 13232: data <= 'd2; 13233: data <= 'd2; 13234: data <= 'd5; 13235: data <= 'd5; 13236: data <= 'd4; 13237: data <= 'd2; 13238: data <= 'd0; 13239: data <= 'd0; 13240: data <= 'd0; 13241: data <= 'd0; 13242: data <= 'd0; 13243: data <= 'd0; 13244: data <= 'd0; 13245: data <= 'd0; 13246: data <= 'd0; 13247: data <= 'd0; 13248: data <= 'd0; 13249: data <= 'd0; 13250: data <= 'd0; 13251: data <= 'd0; 13252: data <= 'd0; 13253: data <= 'd0; 13254: data <= 'd0; 13255: data <= 'd0; 13256: data <= 'd0; 13257: data <= 'd0; 13258: data <= 'd0; 13259: data <= 'd2; 13260: data <= 'd4; 13261: data <= 'd7; 13262: data <= 'd2; 13263: data <= 'd0; 13264: data <= 'd0; 13265: data <= 'd0; 13266: data <= 'd2; 13267: data <= 'd4; 13268: data <= 'd4; 13269: data <= 'd2; 13270: data <= 'd0; 13271: data <= 'd0; 13272: data <= 'd0; 13273: data <= 'd0; 13274: data <= 'd0; 13275: data <= 'd0; 13276: data <= 'd0; 13277: data <= 'd0; 13278: data <= 'd0; 13279: data <= 'd0; 13280: data <= 'd0; 13281: data <= 'd0; 13282: data <= 'd0; 13283: data <= 'd0; 13284: data <= 'd0; 13285: data <= 'd0; 13286: data <= 'd0; 13287: data <= 'd0; 13288: data <= 'd0; 13289: data <= 'd0; 13290: data <= 'd0; 13291: data <= 'd2; 13292: data <= 'd2; 13293: data <= 'd2; 13294: data <= 'd0; 13295: data <= 'd0; 13296: data <= 'd0; 13297: data <= 'd0; 13298: data <= 'd2; 13299: data <= 'd2; 13300: data <= 'd2; 13301: data <= 'd0; 13302: data <= 'd0; 13303: data <= 'd0; 13304: data <= 'd0; 13305: data <= 'd0; 13306: data <= 'd0; 13307: data <= 'd0; 13308: data <= 'd0; 13309: data <= 'd0; 13310: data <= 'd0; 13311: data <= 'd0; 13312: data <= 'd0; 13313: data <= 'd0; 13314: data <= 'd0; 13315: data <= 'd0; 13316: data <= 'd0; 13317: data <= 'd0; 13318: data <= 'd0; 13319: data <= 'd0; 13320: data <= 'd0; 13321: data <= 'd0; 13322: data <= 'd0; 13323: data <= 'd0; 13324: data <= 'd0; 13325: data <= 'd0; 13326: data <= 'd0; 13327: data <= 'd0; 13328: data <= 'd0; 13329: data <= 'd0; 13330: data <= 'd0; 13331: data <= 'd0; 13332: data <= 'd0; 13333: data <= 'd0; 13334: data <= 'd0; 13335: data <= 'd0; 13336: data <= 'd0; 13337: data <= 'd0; 13338: data <= 'd0; 13339: data <= 'd0; 13340: data <= 'd0; 13341: data <= 'd0; 13342: data <= 'd0; 13343: data <= 'd0; 13344: data <= 'd0; 13345: data <= 'd0; 13346: data <= 'd0; 13347: data <= 'd0; 13348: data <= 'd0; 13349: data <= 'd0; 13350: data <= 'd0; 13351: data <= 'd0; 13352: data <= 'd0; 13353: data <= 'd0; 13354: data <= 'd0; 13355: data <= 'd0; 13356: data <= 'd0; 13357: data <= 'd0; 13358: data <= 'd0; 13359: data <= 'd0; 13360: data <= 'd0; 13361: data <= 'd0; 13362: data <= 'd0; 13363: data <= 'd0; 13364: data <= 'd0; 13365: data <= 'd0; 13366: data <= 'd0; 13367: data <= 'd0; 13368: data <= 'd0; 13369: data <= 'd0; 13370: data <= 'd0; 13371: data <= 'd0; 13372: data <= 'd0; 13373: data <= 'd0; 13374: data <= 'd0; 13375: data <= 'd0; 13376: data <= 'd0; 13377: data <= 'd0; 13378: data <= 'd0; 13379: data <= 'd0; 13380: data <= 'd0; 13381: data <= 'd0; 13382: data <= 'd0; 13383: data <= 'd0; 13384: data <= 'd0; 13385: data <= 'd0; 13386: data <= 'd0; 13387: data <= 'd0; 13388: data <= 'd0; 13389: data <= 'd0; 13390: data <= 'd0; 13391: data <= 'd0; 13392: data <= 'd0; 13393: data <= 'd0; 13394: data <= 'd0; 13395: data <= 'd0; 13396: data <= 'd0; 13397: data <= 'd0; 13398: data <= 'd0; 13399: data <= 'd0; 13400: data <= 'd0; 13401: data <= 'd0; 13402: data <= 'd0; 13403: data <= 'd0; 13404: data <= 'd0; 13405: data <= 'd0; 13406: data <= 'd0; 13407: data <= 'd0; 13408: data <= 'd0; 13409: data <= 'd0; 13410: data <= 'd0; 13411: data <= 'd0; 13412: data <= 'd0; 13413: data <= 'd0; 13414: data <= 'd0; 13415: data <= 'd0; 13416: data <= 'd0; 13417: data <= 'd0; 13418: data <= 'd0; 13419: data <= 'd0; 13420: data <= 'd0; 13421: data <= 'd0; 13422: data <= 'd0; 13423: data <= 'd0; 13424: data <= 'd0; 13425: data <= 'd0; 13426: data <= 'd0; 13427: data <= 'd0; 13428: data <= 'd0; 13429: data <= 'd0; 13430: data <= 'd0; 13431: data <= 'd0; 13432: data <= 'd0; 13433: data <= 'd0; 13434: data <= 'd0; 13435: data <= 'd0; 13436: data <= 'd0; 13437: data <= 'd0; 13438: data <= 'd0; 13439: data <= 'd0; 13440: data <= 'd0; 13441: data <= 'd0; 13442: data <= 'd0; 13443: data <= 'd0; 13444: data <= 'd0; 13445: data <= 'd0; 13446: data <= 'd0; 13447: data <= 'd0; 13448: data <= 'd0; 13449: data <= 'd0; 13450: data <= 'd0; 13451: data <= 'd0; 13452: data <= 'd0; 13453: data <= 'd0; 13454: data <= 'd0; 13455: data <= 'd0; 13456: data <= 'd0; 13457: data <= 'd0; 13458: data <= 'd0; 13459: data <= 'd0; 13460: data <= 'd0; 13461: data <= 'd0; 13462: data <= 'd0; 13463: data <= 'd0; 13464: data <= 'd0; 13465: data <= 'd0; 13466: data <= 'd0; 13467: data <= 'd0; 13468: data <= 'd0; 13469: data <= 'd0; 13470: data <= 'd0; 13471: data <= 'd0; 13472: data <= 'd0; 13473: data <= 'd0; 13474: data <= 'd0; 13475: data <= 'd0; 13476: data <= 'd0; 13477: data <= 'd0; 13478: data <= 'd0; 13479: data <= 'd0; 13480: data <= 'd0; 13481: data <= 'd0; 13482: data <= 'd0; 13483: data <= 'd0; 13484: data <= 'd0; 13485: data <= 'd0; 13486: data <= 'd0; 13487: data <= 'd0; 13488: data <= 'd0; 13489: data <= 'd0; 13490: data <= 'd0; 13491: data <= 'd0; 13492: data <= 'd0; 13493: data <= 'd0; 13494: data <= 'd0; 13495: data <= 'd0; 13496: data <= 'd0; 13497: data <= 'd0; 13498: data <= 'd0; 13499: data <= 'd0; 13500: data <= 'd0; 13501: data <= 'd0; 13502: data <= 'd0; 13503: data <= 'd0; 13504: data <= 'd0; 13505: data <= 'd0; 13506: data <= 'd0; 13507: data <= 'd0; 13508: data <= 'd0; 13509: data <= 'd0; 13510: data <= 'd0; 13511: data <= 'd0; 13512: data <= 'd0; 13513: data <= 'd0; 13514: data <= 'd0; 13515: data <= 'd0; 13516: data <= 'd0; 13517: data <= 'd0; 13518: data <= 'd0; 13519: data <= 'd0; 13520: data <= 'd0; 13521: data <= 'd0; 13522: data <= 'd0; 13523: data <= 'd0; 13524: data <= 'd0; 13525: data <= 'd0; 13526: data <= 'd0; 13527: data <= 'd0; 13528: data <= 'd0; 13529: data <= 'd0; 13530: data <= 'd0; 13531: data <= 'd0; 13532: data <= 'd0; 13533: data <= 'd0; 13534: data <= 'd0; 13535: data <= 'd0; 13536: data <= 'd0; 13537: data <= 'd0; 13538: data <= 'd0; 13539: data <= 'd0; 13540: data <= 'd0; 13541: data <= 'd0; 13542: data <= 'd0; 13543: data <= 'd0; 13544: data <= 'd0; 13545: data <= 'd0; 13546: data <= 'd0; 13547: data <= 'd0; 13548: data <= 'd0; 13549: data <= 'd0; 13550: data <= 'd0; 13551: data <= 'd0; 13552: data <= 'd0; 13553: data <= 'd0; 13554: data <= 'd0; 13555: data <= 'd0; 13556: data <= 'd0; 13557: data <= 'd0; 13558: data <= 'd0; 13559: data <= 'd0; 13560: data <= 'd0; 13561: data <= 'd0; 13562: data <= 'd0; 13563: data <= 'd0; 13564: data <= 'd0; 13565: data <= 'd0; 13566: data <= 'd0; 13567: data <= 'd0; 13568: data <= 'd0; 13569: data <= 'd0; 13570: data <= 'd0; 13571: data <= 'd0; 13572: data <= 'd0; 13573: data <= 'd0; 13574: data <= 'd0; 13575: data <= 'd0; 13576: data <= 'd0; 13577: data <= 'd0; 13578: data <= 'd0; 13579: data <= 'd0; 13580: data <= 'd0; 13581: data <= 'd0; 13582: data <= 'd0; 13583: data <= 'd0; 13584: data <= 'd0; 13585: data <= 'd0; 13586: data <= 'd0; 13587: data <= 'd0; 13588: data <= 'd0; 13589: data <= 'd0; 13590: data <= 'd0; 13591: data <= 'd0; 13592: data <= 'd0; 13593: data <= 'd0; 13594: data <= 'd0; 13595: data <= 'd0; 13596: data <= 'd0; 13597: data <= 'd0; 13598: data <= 'd0; 13599: data <= 'd0; 13600: data <= 'd0; 13601: data <= 'd0; 13602: data <= 'd0; 13603: data <= 'd0; 13604: data <= 'd0; 13605: data <= 'd0; 13606: data <= 'd0; 13607: data <= 'd0; 13608: data <= 'd0; 13609: data <= 'd0; 13610: data <= 'd0; 13611: data <= 'd0; 13612: data <= 'd0; 13613: data <= 'd2; 13614: data <= 'd2; 13615: data <= 'd2; 13616: data <= 'd2; 13617: data <= 'd2; 13618: data <= 'd2; 13619: data <= 'd0; 13620: data <= 'd0; 13621: data <= 'd0; 13622: data <= 'd0; 13623: data <= 'd0; 13624: data <= 'd0; 13625: data <= 'd0; 13626: data <= 'd0; 13627: data <= 'd0; 13628: data <= 'd0; 13629: data <= 'd0; 13630: data <= 'd0; 13631: data <= 'd0; 13632: data <= 'd0; 13633: data <= 'd0; 13634: data <= 'd0; 13635: data <= 'd0; 13636: data <= 'd0; 13637: data <= 'd0; 13638: data <= 'd0; 13639: data <= 'd0; 13640: data <= 'd0; 13641: data <= 'd0; 13642: data <= 'd0; 13643: data <= 'd2; 13644: data <= 'd2; 13645: data <= 'd6; 13646: data <= 'd6; 13647: data <= 'd6; 13648: data <= 'd6; 13649: data <= 'd6; 13650: data <= 'd6; 13651: data <= 'd2; 13652: data <= 'd2; 13653: data <= 'd0; 13654: data <= 'd0; 13655: data <= 'd0; 13656: data <= 'd0; 13657: data <= 'd0; 13658: data <= 'd0; 13659: data <= 'd0; 13660: data <= 'd0; 13661: data <= 'd0; 13662: data <= 'd0; 13663: data <= 'd0; 13664: data <= 'd0; 13665: data <= 'd0; 13666: data <= 'd0; 13667: data <= 'd0; 13668: data <= 'd0; 13669: data <= 'd0; 13670: data <= 'd0; 13671: data <= 'd0; 13672: data <= 'd0; 13673: data <= 'd0; 13674: data <= 'd2; 13675: data <= 'd1; 13676: data <= 'd3; 13677: data <= 'd6; 13678: data <= 'd6; 13679: data <= 'd6; 13680: data <= 'd6; 13681: data <= 'd6; 13682: data <= 'd6; 13683: data <= 'd6; 13684: data <= 'd3; 13685: data <= 'd2; 13686: data <= 'd0; 13687: data <= 'd0; 13688: data <= 'd0; 13689: data <= 'd0; 13690: data <= 'd0; 13691: data <= 'd0; 13692: data <= 'd0; 13693: data <= 'd0; 13694: data <= 'd0; 13695: data <= 'd0; 13696: data <= 'd0; 13697: data <= 'd0; 13698: data <= 'd0; 13699: data <= 'd0; 13700: data <= 'd0; 13701: data <= 'd0; 13702: data <= 'd0; 13703: data <= 'd0; 13704: data <= 'd0; 13705: data <= 'd2; 13706: data <= 'd1; 13707: data <= 'd1; 13708: data <= 'd1; 13709: data <= 'd3; 13710: data <= 'd6; 13711: data <= 'd6; 13712: data <= 'd6; 13713: data <= 'd6; 13714: data <= 'd6; 13715: data <= 'd3; 13716: data <= 'd1; 13717: data <= 'd1; 13718: data <= 'd2; 13719: data <= 'd0; 13720: data <= 'd0; 13721: data <= 'd0; 13722: data <= 'd0; 13723: data <= 'd0; 13724: data <= 'd0; 13725: data <= 'd0; 13726: data <= 'd0; 13727: data <= 'd0; 13728: data <= 'd0; 13729: data <= 'd0; 13730: data <= 'd0; 13731: data <= 'd0; 13732: data <= 'd0; 13733: data <= 'd0; 13734: data <= 'd0; 13735: data <= 'd0; 13736: data <= 'd0; 13737: data <= 'd2; 13738: data <= 'd1; 13739: data <= 'd1; 13740: data <= 'd5; 13741: data <= 'd5; 13742: data <= 'd5; 13743: data <= 'd1; 13744: data <= 'd1; 13745: data <= 'd1; 13746: data <= 'd1; 13747: data <= 'd1; 13748: data <= 'd5; 13749: data <= 'd5; 13750: data <= 'd2; 13751: data <= 'd0; 13752: data <= 'd0; 13753: data <= 'd0; 13754: data <= 'd0; 13755: data <= 'd0; 13756: data <= 'd0; 13757: data <= 'd0; 13758: data <= 'd0; 13759: data <= 'd0; 13760: data <= 'd0; 13761: data <= 'd0; 13762: data <= 'd0; 13763: data <= 'd0; 13764: data <= 'd0; 13765: data <= 'd0; 13766: data <= 'd0; 13767: data <= 'd0; 13768: data <= 'd2; 13769: data <= 'd1; 13770: data <= 'd5; 13771: data <= 'd5; 13772: data <= 'd3; 13773: data <= 'd6; 13774: data <= 'd6; 13775: data <= 'd6; 13776: data <= 'd6; 13777: data <= 'd6; 13778: data <= 'd6; 13779: data <= 'd6; 13780: data <= 'd6; 13781: data <= 'd3; 13782: data <= 'd5; 13783: data <= 'd2; 13784: data <= 'd0; 13785: data <= 'd0; 13786: data <= 'd0; 13787: data <= 'd0; 13788: data <= 'd0; 13789: data <= 'd0; 13790: data <= 'd0; 13791: data <= 'd0; 13792: data <= 'd0; 13793: data <= 'd0; 13794: data <= 'd0; 13795: data <= 'd0; 13796: data <= 'd0; 13797: data <= 'd0; 13798: data <= 'd0; 13799: data <= 'd0; 13800: data <= 'd2; 13801: data <= 'd5; 13802: data <= 'd3; 13803: data <= 'd6; 13804: data <= 'd3; 13805: data <= 'd1; 13806: data <= 'd1; 13807: data <= 'd1; 13808: data <= 'd1; 13809: data <= 'd1; 13810: data <= 'd1; 13811: data <= 'd1; 13812: data <= 'd1; 13813: data <= 'd1; 13814: data <= 'd3; 13815: data <= 'd2; 13816: data <= 'd0; 13817: data <= 'd0; 13818: data <= 'd0; 13819: data <= 'd0; 13820: data <= 'd0; 13821: data <= 'd0; 13822: data <= 'd0; 13823: data <= 'd0; 13824: data <= 'd0; 13825: data <= 'd0; 13826: data <= 'd0; 13827: data <= 'd0; 13828: data <= 'd0; 13829: data <= 'd0; 13830: data <= 'd0; 13831: data <= 'd0; 13832: data <= 'd2; 13833: data <= 'd5; 13834: data <= 'd3; 13835: data <= 'd1; 13836: data <= 'd1; 13837: data <= 'd1; 13838: data <= 'd5; 13839: data <= 'd5; 13840: data <= 'd5; 13841: data <= 'd5; 13842: data <= 'd5; 13843: data <= 'd5; 13844: data <= 'd5; 13845: data <= 'd1; 13846: data <= 'd1; 13847: data <= 'd2; 13848: data <= 'd0; 13849: data <= 'd0; 13850: data <= 'd0; 13851: data <= 'd0; 13852: data <= 'd0; 13853: data <= 'd0; 13854: data <= 'd0; 13855: data <= 'd0; 13856: data <= 'd0; 13857: data <= 'd0; 13858: data <= 'd0; 13859: data <= 'd0; 13860: data <= 'd0; 13861: data <= 'd0; 13862: data <= 'd0; 13863: data <= 'd0; 13864: data <= 'd2; 13865: data <= 'd6; 13866: data <= 'd1; 13867: data <= 'd5; 13868: data <= 'd2; 13869: data <= 'd2; 13870: data <= 'd2; 13871: data <= 'd2; 13872: data <= 'd2; 13873: data <= 'd2; 13874: data <= 'd2; 13875: data <= 'd2; 13876: data <= 'd2; 13877: data <= 'd2; 13878: data <= 'd5; 13879: data <= 'd2; 13880: data <= 'd0; 13881: data <= 'd0; 13882: data <= 'd0; 13883: data <= 'd0; 13884: data <= 'd0; 13885: data <= 'd0; 13886: data <= 'd0; 13887: data <= 'd0; 13888: data <= 'd0; 13889: data <= 'd0; 13890: data <= 'd0; 13891: data <= 'd0; 13892: data <= 'd0; 13893: data <= 'd0; 13894: data <= 'd2; 13895: data <= 'd2; 13896: data <= 'd5; 13897: data <= 'd6; 13898: data <= 'd5; 13899: data <= 'd2; 13900: data <= 'd8; 13901: data <= 'd8; 13902: data <= 'd8; 13903: data <= 'd8; 13904: data <= 'd8; 13905: data <= 'd9; 13906: data <= 'd9; 13907: data <= 'd8; 13908: data <= 'd8; 13909: data <= 'd8; 13910: data <= 'd2; 13911: data <= 'd2; 13912: data <= 'd0; 13913: data <= 'd0; 13914: data <= 'd0; 13915: data <= 'd0; 13916: data <= 'd0; 13917: data <= 'd0; 13918: data <= 'd0; 13919: data <= 'd0; 13920: data <= 'd0; 13921: data <= 'd0; 13922: data <= 'd0; 13923: data <= 'd0; 13924: data <= 'd0; 13925: data <= 'd0; 13926: data <= 'd2; 13927: data <= 'd3; 13928: data <= 'd6; 13929: data <= 'd3; 13930: data <= 'd2; 13931: data <= 'd8; 13932: data <= 'd8; 13933: data <= 'd9; 13934: data <= 'd9; 13935: data <= 'd10; 13936: data <= 'd2; 13937: data <= 'd9; 13938: data <= 'd11; 13939: data <= 'd10; 13940: data <= 'd2; 13941: data <= 'd9; 13942: data <= 'd2; 13943: data <= 'd2; 13944: data <= 'd0; 13945: data <= 'd0; 13946: data <= 'd0; 13947: data <= 'd0; 13948: data <= 'd0; 13949: data <= 'd0; 13950: data <= 'd0; 13951: data <= 'd0; 13952: data <= 'd0; 13953: data <= 'd0; 13954: data <= 'd0; 13955: data <= 'd0; 13956: data <= 'd0; 13957: data <= 'd0; 13958: data <= 'd2; 13959: data <= 'd1; 13960: data <= 'd3; 13961: data <= 'd1; 13962: data <= 'd2; 13963: data <= 'd10; 13964: data <= 'd10; 13965: data <= 'd9; 13966: data <= 'd10; 13967: data <= 'd10; 13968: data <= 'd11; 13969: data <= 'd10; 13970: data <= 'd11; 13971: data <= 'd11; 13972: data <= 'd10; 13973: data <= 'd10; 13974: data <= 'd2; 13975: data <= 'd0; 13976: data <= 'd0; 13977: data <= 'd0; 13978: data <= 'd0; 13979: data <= 'd0; 13980: data <= 'd0; 13981: data <= 'd0; 13982: data <= 'd0; 13983: data <= 'd0; 13984: data <= 'd0; 13985: data <= 'd0; 13986: data <= 'd0; 13987: data <= 'd0; 13988: data <= 'd0; 13989: data <= 'd0; 13990: data <= 'd0; 13991: data <= 'd2; 13992: data <= 'd1; 13993: data <= 'd5; 13994: data <= 'd2; 13995: data <= 'd8; 13996: data <= 'd9; 13997: data <= 'd9; 13998: data <= 'd10; 13999: data <= 'd10; 14000: data <= 'd10; 14001: data <= 'd10; 14002: data <= 'd8; 14003: data <= 'd8; 14004: data <= 'd10; 14005: data <= 'd9; 14006: data <= 'd2; 14007: data <= 'd0; 14008: data <= 'd0; 14009: data <= 'd0; 14010: data <= 'd0; 14011: data <= 'd0; 14012: data <= 'd0; 14013: data <= 'd0; 14014: data <= 'd0; 14015: data <= 'd0; 14016: data <= 'd0; 14017: data <= 'd0; 14018: data <= 'd0; 14019: data <= 'd0; 14020: data <= 'd0; 14021: data <= 'd0; 14022: data <= 'd0; 14023: data <= 'd0; 14024: data <= 'd2; 14025: data <= 'd2; 14026: data <= 'd2; 14027: data <= 'd8; 14028: data <= 'd8; 14029: data <= 'd9; 14030: data <= 'd9; 14031: data <= 'd10; 14032: data <= 'd10; 14033: data <= 'd10; 14034: data <= 'd9; 14035: data <= 'd9; 14036: data <= 'd10; 14037: data <= 'd9; 14038: data <= 'd2; 14039: data <= 'd0; 14040: data <= 'd0; 14041: data <= 'd0; 14042: data <= 'd0; 14043: data <= 'd0; 14044: data <= 'd0; 14045: data <= 'd0; 14046: data <= 'd0; 14047: data <= 'd0; 14048: data <= 'd0; 14049: data <= 'd0; 14050: data <= 'd0; 14051: data <= 'd0; 14052: data <= 'd0; 14053: data <= 'd0; 14054: data <= 'd0; 14055: data <= 'd0; 14056: data <= 'd0; 14057: data <= 'd0; 14058: data <= 'd0; 14059: data <= 'd2; 14060: data <= 'd5; 14061: data <= 'd5; 14062: data <= 'd8; 14063: data <= 'd9; 14064: data <= 'd9; 14065: data <= 'd9; 14066: data <= 'd9; 14067: data <= 'd9; 14068: data <= 'd9; 14069: data <= 'd5; 14070: data <= 'd2; 14071: data <= 'd0; 14072: data <= 'd0; 14073: data <= 'd0; 14074: data <= 'd0; 14075: data <= 'd0; 14076: data <= 'd0; 14077: data <= 'd0; 14078: data <= 'd0; 14079: data <= 'd0; 14080: data <= 'd0; 14081: data <= 'd0; 14082: data <= 'd0; 14083: data <= 'd0; 14084: data <= 'd0; 14085: data <= 'd0; 14086: data <= 'd0; 14087: data <= 'd0; 14088: data <= 'd0; 14089: data <= 'd0; 14090: data <= 'd0; 14091: data <= 'd2; 14092: data <= 'd1; 14093: data <= 'd1; 14094: data <= 'd3; 14095: data <= 'd3; 14096: data <= 'd5; 14097: data <= 'd5; 14098: data <= 'd3; 14099: data <= 'd3; 14100: data <= 'd1; 14101: data <= 'd2; 14102: data <= 'd0; 14103: data <= 'd0; 14104: data <= 'd0; 14105: data <= 'd0; 14106: data <= 'd0; 14107: data <= 'd0; 14108: data <= 'd0; 14109: data <= 'd0; 14110: data <= 'd0; 14111: data <= 'd0; 14112: data <= 'd0; 14113: data <= 'd0; 14114: data <= 'd0; 14115: data <= 'd0; 14116: data <= 'd0; 14117: data <= 'd0; 14118: data <= 'd0; 14119: data <= 'd0; 14120: data <= 'd0; 14121: data <= 'd0; 14122: data <= 'd0; 14123: data <= 'd2; 14124: data <= 'd7; 14125: data <= 'd1; 14126: data <= 'd5; 14127: data <= 'd5; 14128: data <= 'd2; 14129: data <= 'd1; 14130: data <= 'd3; 14131: data <= 'd3; 14132: data <= 'd1; 14133: data <= 'd2; 14134: data <= 'd0; 14135: data <= 'd0; 14136: data <= 'd0; 14137: data <= 'd0; 14138: data <= 'd0; 14139: data <= 'd0; 14140: data <= 'd0; 14141: data <= 'd0; 14142: data <= 'd0; 14143: data <= 'd0; 14144: data <= 'd0; 14145: data <= 'd0; 14146: data <= 'd0; 14147: data <= 'd0; 14148: data <= 'd0; 14149: data <= 'd0; 14150: data <= 'd0; 14151: data <= 'd0; 14152: data <= 'd0; 14153: data <= 'd0; 14154: data <= 'd0; 14155: data <= 'd2; 14156: data <= 'd2; 14157: data <= 'd7; 14158: data <= 'd10; 14159: data <= 'd10; 14160: data <= 'd10; 14161: data <= 'd2; 14162: data <= 'd3; 14163: data <= 'd1; 14164: data <= 'd1; 14165: data <= 'd2; 14166: data <= 'd0; 14167: data <= 'd0; 14168: data <= 'd0; 14169: data <= 'd0; 14170: data <= 'd0; 14171: data <= 'd0; 14172: data <= 'd0; 14173: data <= 'd0; 14174: data <= 'd0; 14175: data <= 'd0; 14176: data <= 'd0; 14177: data <= 'd0; 14178: data <= 'd0; 14179: data <= 'd0; 14180: data <= 'd0; 14181: data <= 'd0; 14182: data <= 'd0; 14183: data <= 'd0; 14184: data <= 'd0; 14185: data <= 'd0; 14186: data <= 'd0; 14187: data <= 'd2; 14188: data <= 'd4; 14189: data <= 'd2; 14190: data <= 'd9; 14191: data <= 'd10; 14192: data <= 'd9; 14193: data <= 'd2; 14194: data <= 'd2; 14195: data <= 'd2; 14196: data <= 'd2; 14197: data <= 'd2; 14198: data <= 'd0; 14199: data <= 'd0; 14200: data <= 'd0; 14201: data <= 'd0; 14202: data <= 'd0; 14203: data <= 'd0; 14204: data <= 'd0; 14205: data <= 'd0; 14206: data <= 'd0; 14207: data <= 'd0; 14208: data <= 'd0; 14209: data <= 'd0; 14210: data <= 'd0; 14211: data <= 'd0; 14212: data <= 'd0; 14213: data <= 'd0; 14214: data <= 'd0; 14215: data <= 'd0; 14216: data <= 'd0; 14217: data <= 'd0; 14218: data <= 'd0; 14219: data <= 'd2; 14220: data <= 'd4; 14221: data <= 'd4; 14222: data <= 'd2; 14223: data <= 'd2; 14224: data <= 'd2; 14225: data <= 'd3; 14226: data <= 'd3; 14227: data <= 'd3; 14228: data <= 'd5; 14229: data <= 'd0; 14230: data <= 'd0; 14231: data <= 'd0; 14232: data <= 'd0; 14233: data <= 'd0; 14234: data <= 'd0; 14235: data <= 'd0; 14236: data <= 'd0; 14237: data <= 'd0; 14238: data <= 'd0; 14239: data <= 'd0; 14240: data <= 'd0; 14241: data <= 'd0; 14242: data <= 'd0; 14243: data <= 'd0; 14244: data <= 'd0; 14245: data <= 'd0; 14246: data <= 'd0; 14247: data <= 'd0; 14248: data <= 'd0; 14249: data <= 'd0; 14250: data <= 'd0; 14251: data <= 'd2; 14252: data <= 'd4; 14253: data <= 'd7; 14254: data <= 'd7; 14255: data <= 'd2; 14256: data <= 'd2; 14257: data <= 'd5; 14258: data <= 'd5; 14259: data <= 'd4; 14260: data <= 'd2; 14261: data <= 'd0; 14262: data <= 'd0; 14263: data <= 'd0; 14264: data <= 'd0; 14265: data <= 'd0; 14266: data <= 'd0; 14267: data <= 'd0; 14268: data <= 'd0; 14269: data <= 'd0; 14270: data <= 'd0; 14271: data <= 'd0; 14272: data <= 'd0; 14273: data <= 'd0; 14274: data <= 'd0; 14275: data <= 'd0; 14276: data <= 'd0; 14277: data <= 'd0; 14278: data <= 'd0; 14279: data <= 'd0; 14280: data <= 'd0; 14281: data <= 'd0; 14282: data <= 'd0; 14283: data <= 'd2; 14284: data <= 'd4; 14285: data <= 'd7; 14286: data <= 'd2; 14287: data <= 'd0; 14288: data <= 'd2; 14289: data <= 'd4; 14290: data <= 'd4; 14291: data <= 'd2; 14292: data <= 'd0; 14293: data <= 'd0; 14294: data <= 'd0; 14295: data <= 'd0; 14296: data <= 'd0; 14297: data <= 'd0; 14298: data <= 'd0; 14299: data <= 'd0; 14300: data <= 'd0; 14301: data <= 'd0; 14302: data <= 'd0; 14303: data <= 'd0; 14304: data <= 'd0; 14305: data <= 'd0; 14306: data <= 'd0; 14307: data <= 'd0; 14308: data <= 'd0; 14309: data <= 'd0; 14310: data <= 'd0; 14311: data <= 'd0; 14312: data <= 'd0; 14313: data <= 'd0; 14314: data <= 'd0; 14315: data <= 'd2; 14316: data <= 'd2; 14317: data <= 'd2; 14318: data <= 'd0; 14319: data <= 'd0; 14320: data <= 'd2; 14321: data <= 'd2; 14322: data <= 'd2; 14323: data <= 'd0; 14324: data <= 'd0; 14325: data <= 'd0; 14326: data <= 'd0; 14327: data <= 'd0; 14328: data <= 'd0; 14329: data <= 'd0; 14330: data <= 'd0; 14331: data <= 'd0; 14332: data <= 'd0; 14333: data <= 'd0; 14334: data <= 'd0; 14335: data <= 'd0; 14336: data <= 'd0; 14337: data <= 'd0; 14338: data <= 'd0; 14339: data <= 'd0; 14340: data <= 'd0; 14341: data <= 'd0; 14342: data <= 'd0; 14343: data <= 'd0; 14344: data <= 'd0; 14345: data <= 'd0; 14346: data <= 'd0; 14347: data <= 'd0; 14348: data <= 'd0; 14349: data <= 'd0; 14350: data <= 'd0; 14351: data <= 'd0; 14352: data <= 'd0; 14353: data <= 'd0; 14354: data <= 'd0; 14355: data <= 'd0; 14356: data <= 'd0; 14357: data <= 'd0; 14358: data <= 'd0; 14359: data <= 'd0; 14360: data <= 'd0; 14361: data <= 'd0; 14362: data <= 'd0; 14363: data <= 'd0; 14364: data <= 'd0; 14365: data <= 'd0; 14366: data <= 'd0; 14367: data <= 'd0; 14368: data <= 'd0; 14369: data <= 'd0; 14370: data <= 'd0; 14371: data <= 'd0; 14372: data <= 'd0; 14373: data <= 'd0; 14374: data <= 'd0; 14375: data <= 'd0; 14376: data <= 'd0; 14377: data <= 'd0; 14378: data <= 'd0; 14379: data <= 'd0; 14380: data <= 'd0; 14381: data <= 'd0; 14382: data <= 'd0; 14383: data <= 'd0; 14384: data <= 'd0; 14385: data <= 'd0; 14386: data <= 'd0; 14387: data <= 'd0; 14388: data <= 'd0; 14389: data <= 'd0; 14390: data <= 'd0; 14391: data <= 'd0; 14392: data <= 'd0; 14393: data <= 'd0; 14394: data <= 'd0; 14395: data <= 'd0; 14396: data <= 'd0; 14397: data <= 'd0; 14398: data <= 'd0; 14399: data <= 'd0; 14400: data <= 'd0; 14401: data <= 'd0; 14402: data <= 'd0; 14403: data <= 'd0; 14404: data <= 'd0; 14405: data <= 'd0; 14406: data <= 'd0; 14407: data <= 'd0; 14408: data <= 'd0; 14409: data <= 'd0; 14410: data <= 'd0; 14411: data <= 'd0; 14412: data <= 'd0; 14413: data <= 'd0; 14414: data <= 'd0; 14415: data <= 'd0; 14416: data <= 'd0; 14417: data <= 'd0; 14418: data <= 'd0; 14419: data <= 'd0; 14420: data <= 'd0; 14421: data <= 'd0; 14422: data <= 'd0; 14423: data <= 'd0; 14424: data <= 'd0; 14425: data <= 'd0; 14426: data <= 'd0; 14427: data <= 'd0; 14428: data <= 'd0; 14429: data <= 'd0; 14430: data <= 'd0; 14431: data <= 'd0; 14432: data <= 'd0; 14433: data <= 'd0; 14434: data <= 'd0; 14435: data <= 'd0; 14436: data <= 'd0; 14437: data <= 'd0; 14438: data <= 'd0; 14439: data <= 'd0; 14440: data <= 'd0; 14441: data <= 'd0; 14442: data <= 'd0; 14443: data <= 'd0; 14444: data <= 'd0; 14445: data <= 'd0; 14446: data <= 'd0; 14447: data <= 'd0; 14448: data <= 'd0; 14449: data <= 'd0; 14450: data <= 'd0; 14451: data <= 'd0; 14452: data <= 'd0; 14453: data <= 'd0; 14454: data <= 'd0; 14455: data <= 'd0; 14456: data <= 'd0; 14457: data <= 'd0; 14458: data <= 'd0; 14459: data <= 'd0; 14460: data <= 'd0; 14461: data <= 'd0; 14462: data <= 'd0; 14463: data <= 'd0; 14464: data <= 'd0; 14465: data <= 'd0; 14466: data <= 'd0; 14467: data <= 'd0; 14468: data <= 'd0; 14469: data <= 'd0; 14470: data <= 'd0; 14471: data <= 'd0; 14472: data <= 'd0; 14473: data <= 'd0; 14474: data <= 'd0; 14475: data <= 'd0; 14476: data <= 'd0; 14477: data <= 'd0; 14478: data <= 'd0; 14479: data <= 'd0; 14480: data <= 'd0; 14481: data <= 'd0; 14482: data <= 'd0; 14483: data <= 'd0; 14484: data <= 'd0; 14485: data <= 'd0; 14486: data <= 'd0; 14487: data <= 'd0; 14488: data <= 'd0; 14489: data <= 'd0; 14490: data <= 'd0; 14491: data <= 'd0; 14492: data <= 'd0; 14493: data <= 'd0; 14494: data <= 'd0; 14495: data <= 'd0; 14496: data <= 'd0; 14497: data <= 'd0; 14498: data <= 'd0; 14499: data <= 'd0; 14500: data <= 'd0; 14501: data <= 'd0; 14502: data <= 'd0; 14503: data <= 'd0; 14504: data <= 'd0; 14505: data <= 'd0; 14506: data <= 'd0; 14507: data <= 'd0; 14508: data <= 'd0; 14509: data <= 'd0; 14510: data <= 'd0; 14511: data <= 'd0; 14512: data <= 'd0; 14513: data <= 'd0; 14514: data <= 'd0; 14515: data <= 'd0; 14516: data <= 'd0; 14517: data <= 'd0; 14518: data <= 'd0; 14519: data <= 'd0; 14520: data <= 'd0; 14521: data <= 'd0; 14522: data <= 'd0; 14523: data <= 'd0; 14524: data <= 'd0; 14525: data <= 'd0; 14526: data <= 'd0; 14527: data <= 'd0; 14528: data <= 'd0; 14529: data <= 'd0; 14530: data <= 'd0; 14531: data <= 'd0; 14532: data <= 'd0; 14533: data <= 'd0; 14534: data <= 'd0; 14535: data <= 'd0; 14536: data <= 'd0; 14537: data <= 'd0; 14538: data <= 'd0; 14539: data <= 'd0; 14540: data <= 'd0; 14541: data <= 'd0; 14542: data <= 'd0; 14543: data <= 'd0; 14544: data <= 'd0; 14545: data <= 'd0; 14546: data <= 'd0; 14547: data <= 'd0; 14548: data <= 'd0; 14549: data <= 'd0; 14550: data <= 'd0; 14551: data <= 'd0; 14552: data <= 'd0; 14553: data <= 'd0; 14554: data <= 'd0; 14555: data <= 'd0; 14556: data <= 'd0; 14557: data <= 'd0; 14558: data <= 'd0; 14559: data <= 'd0; 14560: data <= 'd0; 14561: data <= 'd0; 14562: data <= 'd0; 14563: data <= 'd0; 14564: data <= 'd0; 14565: data <= 'd0; 14566: data <= 'd0; 14567: data <= 'd0; 14568: data <= 'd0; 14569: data <= 'd0; 14570: data <= 'd0; 14571: data <= 'd0; 14572: data <= 'd0; 14573: data <= 'd0; 14574: data <= 'd0; 14575: data <= 'd0; 14576: data <= 'd0; 14577: data <= 'd0; 14578: data <= 'd0; 14579: data <= 'd0; 14580: data <= 'd0; 14581: data <= 'd0; 14582: data <= 'd0; 14583: data <= 'd0; 14584: data <= 'd0; 14585: data <= 'd0; 14586: data <= 'd0; 14587: data <= 'd0; 14588: data <= 'd0; 14589: data <= 'd0; 14590: data <= 'd0; 14591: data <= 'd0; 14592: data <= 'd0; 14593: data <= 'd0; 14594: data <= 'd0; 14595: data <= 'd0; 14596: data <= 'd0; 14597: data <= 'd0; 14598: data <= 'd0; 14599: data <= 'd0; 14600: data <= 'd0; 14601: data <= 'd0; 14602: data <= 'd0; 14603: data <= 'd0; 14604: data <= 'd0; 14605: data <= 'd2; 14606: data <= 'd2; 14607: data <= 'd2; 14608: data <= 'd2; 14609: data <= 'd2; 14610: data <= 'd2; 14611: data <= 'd0; 14612: data <= 'd0; 14613: data <= 'd0; 14614: data <= 'd0; 14615: data <= 'd0; 14616: data <= 'd0; 14617: data <= 'd0; 14618: data <= 'd0; 14619: data <= 'd0; 14620: data <= 'd0; 14621: data <= 'd0; 14622: data <= 'd0; 14623: data <= 'd0; 14624: data <= 'd0; 14625: data <= 'd0; 14626: data <= 'd0; 14627: data <= 'd0; 14628: data <= 'd0; 14629: data <= 'd0; 14630: data <= 'd0; 14631: data <= 'd0; 14632: data <= 'd0; 14633: data <= 'd0; 14634: data <= 'd0; 14635: data <= 'd2; 14636: data <= 'd2; 14637: data <= 'd6; 14638: data <= 'd6; 14639: data <= 'd6; 14640: data <= 'd6; 14641: data <= 'd6; 14642: data <= 'd6; 14643: data <= 'd2; 14644: data <= 'd2; 14645: data <= 'd0; 14646: data <= 'd0; 14647: data <= 'd0; 14648: data <= 'd0; 14649: data <= 'd0; 14650: data <= 'd0; 14651: data <= 'd0; 14652: data <= 'd0; 14653: data <= 'd0; 14654: data <= 'd0; 14655: data <= 'd0; 14656: data <= 'd0; 14657: data <= 'd0; 14658: data <= 'd0; 14659: data <= 'd0; 14660: data <= 'd0; 14661: data <= 'd0; 14662: data <= 'd0; 14663: data <= 'd0; 14664: data <= 'd0; 14665: data <= 'd0; 14666: data <= 'd2; 14667: data <= 'd1; 14668: data <= 'd3; 14669: data <= 'd6; 14670: data <= 'd6; 14671: data <= 'd6; 14672: data <= 'd6; 14673: data <= 'd6; 14674: data <= 'd6; 14675: data <= 'd6; 14676: data <= 'd3; 14677: data <= 'd2; 14678: data <= 'd0; 14679: data <= 'd0; 14680: data <= 'd0; 14681: data <= 'd0; 14682: data <= 'd0; 14683: data <= 'd0; 14684: data <= 'd0; 14685: data <= 'd0; 14686: data <= 'd0; 14687: data <= 'd0; 14688: data <= 'd0; 14689: data <= 'd0; 14690: data <= 'd0; 14691: data <= 'd0; 14692: data <= 'd0; 14693: data <= 'd0; 14694: data <= 'd0; 14695: data <= 'd0; 14696: data <= 'd0; 14697: data <= 'd2; 14698: data <= 'd1; 14699: data <= 'd1; 14700: data <= 'd1; 14701: data <= 'd3; 14702: data <= 'd6; 14703: data <= 'd6; 14704: data <= 'd6; 14705: data <= 'd6; 14706: data <= 'd6; 14707: data <= 'd3; 14708: data <= 'd1; 14709: data <= 'd1; 14710: data <= 'd2; 14711: data <= 'd0; 14712: data <= 'd0; 14713: data <= 'd0; 14714: data <= 'd0; 14715: data <= 'd0; 14716: data <= 'd0; 14717: data <= 'd0; 14718: data <= 'd0; 14719: data <= 'd0; 14720: data <= 'd0; 14721: data <= 'd0; 14722: data <= 'd0; 14723: data <= 'd0; 14724: data <= 'd0; 14725: data <= 'd0; 14726: data <= 'd0; 14727: data <= 'd0; 14728: data <= 'd0; 14729: data <= 'd2; 14730: data <= 'd1; 14731: data <= 'd1; 14732: data <= 'd5; 14733: data <= 'd5; 14734: data <= 'd5; 14735: data <= 'd1; 14736: data <= 'd1; 14737: data <= 'd1; 14738: data <= 'd1; 14739: data <= 'd1; 14740: data <= 'd5; 14741: data <= 'd5; 14742: data <= 'd2; 14743: data <= 'd0; 14744: data <= 'd0; 14745: data <= 'd0; 14746: data <= 'd0; 14747: data <= 'd0; 14748: data <= 'd0; 14749: data <= 'd0; 14750: data <= 'd0; 14751: data <= 'd0; 14752: data <= 'd0; 14753: data <= 'd0; 14754: data <= 'd0; 14755: data <= 'd0; 14756: data <= 'd0; 14757: data <= 'd0; 14758: data <= 'd0; 14759: data <= 'd0; 14760: data <= 'd2; 14761: data <= 'd1; 14762: data <= 'd5; 14763: data <= 'd5; 14764: data <= 'd3; 14765: data <= 'd6; 14766: data <= 'd6; 14767: data <= 'd6; 14768: data <= 'd6; 14769: data <= 'd6; 14770: data <= 'd6; 14771: data <= 'd6; 14772: data <= 'd6; 14773: data <= 'd3; 14774: data <= 'd5; 14775: data <= 'd2; 14776: data <= 'd0; 14777: data <= 'd0; 14778: data <= 'd0; 14779: data <= 'd0; 14780: data <= 'd0; 14781: data <= 'd0; 14782: data <= 'd0; 14783: data <= 'd0; 14784: data <= 'd0; 14785: data <= 'd0; 14786: data <= 'd0; 14787: data <= 'd0; 14788: data <= 'd0; 14789: data <= 'd0; 14790: data <= 'd0; 14791: data <= 'd0; 14792: data <= 'd2; 14793: data <= 'd5; 14794: data <= 'd3; 14795: data <= 'd6; 14796: data <= 'd3; 14797: data <= 'd1; 14798: data <= 'd1; 14799: data <= 'd1; 14800: data <= 'd1; 14801: data <= 'd1; 14802: data <= 'd1; 14803: data <= 'd1; 14804: data <= 'd1; 14805: data <= 'd1; 14806: data <= 'd3; 14807: data <= 'd2; 14808: data <= 'd0; 14809: data <= 'd0; 14810: data <= 'd0; 14811: data <= 'd0; 14812: data <= 'd0; 14813: data <= 'd0; 14814: data <= 'd0; 14815: data <= 'd0; 14816: data <= 'd0; 14817: data <= 'd0; 14818: data <= 'd0; 14819: data <= 'd0; 14820: data <= 'd0; 14821: data <= 'd0; 14822: data <= 'd0; 14823: data <= 'd0; 14824: data <= 'd2; 14825: data <= 'd5; 14826: data <= 'd3; 14827: data <= 'd1; 14828: data <= 'd1; 14829: data <= 'd1; 14830: data <= 'd5; 14831: data <= 'd5; 14832: data <= 'd5; 14833: data <= 'd5; 14834: data <= 'd5; 14835: data <= 'd5; 14836: data <= 'd5; 14837: data <= 'd1; 14838: data <= 'd1; 14839: data <= 'd2; 14840: data <= 'd0; 14841: data <= 'd0; 14842: data <= 'd0; 14843: data <= 'd0; 14844: data <= 'd0; 14845: data <= 'd0; 14846: data <= 'd0; 14847: data <= 'd0; 14848: data <= 'd0; 14849: data <= 'd0; 14850: data <= 'd0; 14851: data <= 'd0; 14852: data <= 'd0; 14853: data <= 'd0; 14854: data <= 'd0; 14855: data <= 'd0; 14856: data <= 'd2; 14857: data <= 'd6; 14858: data <= 'd1; 14859: data <= 'd5; 14860: data <= 'd2; 14861: data <= 'd2; 14862: data <= 'd2; 14863: data <= 'd2; 14864: data <= 'd2; 14865: data <= 'd2; 14866: data <= 'd2; 14867: data <= 'd2; 14868: data <= 'd2; 14869: data <= 'd2; 14870: data <= 'd5; 14871: data <= 'd2; 14872: data <= 'd0; 14873: data <= 'd0; 14874: data <= 'd0; 14875: data <= 'd0; 14876: data <= 'd0; 14877: data <= 'd0; 14878: data <= 'd0; 14879: data <= 'd0; 14880: data <= 'd0; 14881: data <= 'd0; 14882: data <= 'd0; 14883: data <= 'd0; 14884: data <= 'd0; 14885: data <= 'd0; 14886: data <= 'd2; 14887: data <= 'd2; 14888: data <= 'd2; 14889: data <= 'd1; 14890: data <= 'd5; 14891: data <= 'd2; 14892: data <= 'd8; 14893: data <= 'd8; 14894: data <= 'd8; 14895: data <= 'd8; 14896: data <= 'd8; 14897: data <= 'd9; 14898: data <= 'd9; 14899: data <= 'd8; 14900: data <= 'd8; 14901: data <= 'd8; 14902: data <= 'd2; 14903: data <= 'd2; 14904: data <= 'd0; 14905: data <= 'd0; 14906: data <= 'd0; 14907: data <= 'd0; 14908: data <= 'd0; 14909: data <= 'd0; 14910: data <= 'd0; 14911: data <= 'd0; 14912: data <= 'd0; 14913: data <= 'd0; 14914: data <= 'd0; 14915: data <= 'd0; 14916: data <= 'd0; 14917: data <= 'd0; 14918: data <= 'd2; 14919: data <= 'd1; 14920: data <= 'd2; 14921: data <= 'd1; 14922: data <= 'd2; 14923: data <= 'd8; 14924: data <= 'd8; 14925: data <= 'd9; 14926: data <= 'd9; 14927: data <= 'd2; 14928: data <= 'd9; 14929: data <= 'd11; 14930: data <= 'd11; 14931: data <= 'd10; 14932: data <= 'd2; 14933: data <= 'd9; 14934: data <= 'd2; 14935: data <= 'd2; 14936: data <= 'd0; 14937: data <= 'd0; 14938: data <= 'd0; 14939: data <= 'd0; 14940: data <= 'd0; 14941: data <= 'd0; 14942: data <= 'd0; 14943: data <= 'd0; 14944: data <= 'd0; 14945: data <= 'd0; 14946: data <= 'd0; 14947: data <= 'd0; 14948: data <= 'd0; 14949: data <= 'd0; 14950: data <= 'd2; 14951: data <= 'd5; 14952: data <= 'd1; 14953: data <= 'd2; 14954: data <= 'd9; 14955: data <= 'd10; 14956: data <= 'd9; 14957: data <= 'd9; 14958: data <= 'd10; 14959: data <= 'd11; 14960: data <= 'd10; 14961: data <= 'd11; 14962: data <= 'd11; 14963: data <= 'd10; 14964: data <= 'd11; 14965: data <= 'd10; 14966: data <= 'd9; 14967: data <= 'd2; 14968: data <= 'd0; 14969: data <= 'd0; 14970: data <= 'd0; 14971: data <= 'd0; 14972: data <= 'd0; 14973: data <= 'd0; 14974: data <= 'd0; 14975: data <= 'd0; 14976: data <= 'd0; 14977: data <= 'd0; 14978: data <= 'd0; 14979: data <= 'd0; 14980: data <= 'd0; 14981: data <= 'd0; 14982: data <= 'd0; 14983: data <= 'd2; 14984: data <= 'd5; 14985: data <= 'd5; 14986: data <= 'd2; 14987: data <= 'd8; 14988: data <= 'd9; 14989: data <= 'd9; 14990: data <= 'd10; 14991: data <= 'd10; 14992: data <= 'd10; 14993: data <= 'd8; 14994: data <= 'd8; 14995: data <= 'd10; 14996: data <= 'd10; 14997: data <= 'd9; 14998: data <= 'd2; 14999: data <= 'd0; 15000: data <= 'd0; 15001: data <= 'd0; 15002: data <= 'd0; 15003: data <= 'd0; 15004: data <= 'd0; 15005: data <= 'd0; 15006: data <= 'd0; 15007: data <= 'd0; 15008: data <= 'd0; 15009: data <= 'd0; 15010: data <= 'd0; 15011: data <= 'd0; 15012: data <= 'd0; 15013: data <= 'd0; 15014: data <= 'd0; 15015: data <= 'd0; 15016: data <= 'd2; 15017: data <= 'd2; 15018: data <= 'd2; 15019: data <= 'd8; 15020: data <= 'd8; 15021: data <= 'd9; 15022: data <= 'd9; 15023: data <= 'd10; 15024: data <= 'd10; 15025: data <= 'd9; 15026: data <= 'd9; 15027: data <= 'd10; 15028: data <= 'd10; 15029: data <= 'd9; 15030: data <= 'd2; 15031: data <= 'd0; 15032: data <= 'd0; 15033: data <= 'd0; 15034: data <= 'd0; 15035: data <= 'd0; 15036: data <= 'd0; 15037: data <= 'd0; 15038: data <= 'd0; 15039: data <= 'd0; 15040: data <= 'd0; 15041: data <= 'd0; 15042: data <= 'd0; 15043: data <= 'd0; 15044: data <= 'd0; 15045: data <= 'd0; 15046: data <= 'd0; 15047: data <= 'd0; 15048: data <= 'd0; 15049: data <= 'd0; 15050: data <= 'd2; 15051: data <= 'd2; 15052: data <= 'd5; 15053: data <= 'd5; 15054: data <= 'd8; 15055: data <= 'd9; 15056: data <= 'd9; 15057: data <= 'd9; 15058: data <= 'd9; 15059: data <= 'd9; 15060: data <= 'd9; 15061: data <= 'd5; 15062: data <= 'd2; 15063: data <= 'd0; 15064: data <= 'd0; 15065: data <= 'd0; 15066: data <= 'd0; 15067: data <= 'd0; 15068: data <= 'd0; 15069: data <= 'd0; 15070: data <= 'd0; 15071: data <= 'd0; 15072: data <= 'd0; 15073: data <= 'd0; 15074: data <= 'd0; 15075: data <= 'd0; 15076: data <= 'd0; 15077: data <= 'd0; 15078: data <= 'd0; 15079: data <= 'd0; 15080: data <= 'd0; 15081: data <= 'd2; 15082: data <= 'd7; 15083: data <= 'd1; 15084: data <= 'd1; 15085: data <= 'd1; 15086: data <= 'd3; 15087: data <= 'd3; 15088: data <= 'd3; 15089: data <= 'd5; 15090: data <= 'd5; 15091: data <= 'd3; 15092: data <= 'd3; 15093: data <= 'd1; 15094: data <= 'd2; 15095: data <= 'd0; 15096: data <= 'd0; 15097: data <= 'd0; 15098: data <= 'd0; 15099: data <= 'd0; 15100: data <= 'd0; 15101: data <= 'd0; 15102: data <= 'd0; 15103: data <= 'd0; 15104: data <= 'd0; 15105: data <= 'd0; 15106: data <= 'd0; 15107: data <= 'd0; 15108: data <= 'd0; 15109: data <= 'd0; 15110: data <= 'd0; 15111: data <= 'd0; 15112: data <= 'd0; 15113: data <= 'd2; 15114: data <= 'd7; 15115: data <= 'd7; 15116: data <= 'd5; 15117: data <= 'd1; 15118: data <= 'd3; 15119: data <= 'd3; 15120: data <= 'd3; 15121: data <= 'd1; 15122: data <= 'd1; 15123: data <= 'd3; 15124: data <= 'd3; 15125: data <= 'd1; 15126: data <= 'd2; 15127: data <= 'd0; 15128: data <= 'd0; 15129: data <= 'd0; 15130: data <= 'd0; 15131: data <= 'd0; 15132: data <= 'd0; 15133: data <= 'd0; 15134: data <= 'd0; 15135: data <= 'd0; 15136: data <= 'd0; 15137: data <= 'd0; 15138: data <= 'd0; 15139: data <= 'd0; 15140: data <= 'd0; 15141: data <= 'd0; 15142: data <= 'd0; 15143: data <= 'd0; 15144: data <= 'd0; 15145: data <= 'd0; 15146: data <= 'd2; 15147: data <= 'd9; 15148: data <= 'd9; 15149: data <= 'd2; 15150: data <= 'd1; 15151: data <= 'd3; 15152: data <= 'd3; 15153: data <= 'd1; 15154: data <= 'd1; 15155: data <= 'd3; 15156: data <= 'd1; 15157: data <= 'd1; 15158: data <= 'd2; 15159: data <= 'd0; 15160: data <= 'd0; 15161: data <= 'd0; 15162: data <= 'd0; 15163: data <= 'd0; 15164: data <= 'd0; 15165: data <= 'd0; 15166: data <= 'd0; 15167: data <= 'd0; 15168: data <= 'd0; 15169: data <= 'd0; 15170: data <= 'd0; 15171: data <= 'd0; 15172: data <= 'd0; 15173: data <= 'd0; 15174: data <= 'd0; 15175: data <= 'd0; 15176: data <= 'd0; 15177: data <= 'd0; 15178: data <= 'd2; 15179: data <= 'd9; 15180: data <= 'd9; 15181: data <= 'd2; 15182: data <= 'd2; 15183: data <= 'd2; 15184: data <= 'd5; 15185: data <= 'd5; 15186: data <= 'd5; 15187: data <= 'd2; 15188: data <= 'd2; 15189: data <= 'd2; 15190: data <= 'd2; 15191: data <= 'd0; 15192: data <= 'd0; 15193: data <= 'd0; 15194: data <= 'd0; 15195: data <= 'd0; 15196: data <= 'd0; 15197: data <= 'd0; 15198: data <= 'd0; 15199: data <= 'd0; 15200: data <= 'd0; 15201: data <= 'd0; 15202: data <= 'd0; 15203: data <= 'd0; 15204: data <= 'd0; 15205: data <= 'd0; 15206: data <= 'd0; 15207: data <= 'd0; 15208: data <= 'd0; 15209: data <= 'd0; 15210: data <= 'd0; 15211: data <= 'd2; 15212: data <= 'd2; 15213: data <= 'd1; 15214: data <= 'd3; 15215: data <= 'd3; 15216: data <= 'd3; 15217: data <= 'd1; 15218: data <= 'd3; 15219: data <= 'd3; 15220: data <= 'd3; 15221: data <= 'd5; 15222: data <= 'd2; 15223: data <= 'd0; 15224: data <= 'd0; 15225: data <= 'd0; 15226: data <= 'd0; 15227: data <= 'd0; 15228: data <= 'd0; 15229: data <= 'd0; 15230: data <= 'd0; 15231: data <= 'd0; 15232: data <= 'd0; 15233: data <= 'd0; 15234: data <= 'd0; 15235: data <= 'd0; 15236: data <= 'd0; 15237: data <= 'd0; 15238: data <= 'd0; 15239: data <= 'd0; 15240: data <= 'd0; 15241: data <= 'd0; 15242: data <= 'd0; 15243: data <= 'd2; 15244: data <= 'd4; 15245: data <= 'd7; 15246: data <= 'd7; 15247: data <= 'd2; 15248: data <= 'd2; 15249: data <= 'd2; 15250: data <= 'd2; 15251: data <= 'd5; 15252: data <= 'd5; 15253: data <= 'd4; 15254: data <= 'd2; 15255: data <= 'd0; 15256: data <= 'd0; 15257: data <= 'd0; 15258: data <= 'd0; 15259: data <= 'd0; 15260: data <= 'd0; 15261: data <= 'd0; 15262: data <= 'd0; 15263: data <= 'd0; 15264: data <= 'd0; 15265: data <= 'd0; 15266: data <= 'd0; 15267: data <= 'd0; 15268: data <= 'd0; 15269: data <= 'd0; 15270: data <= 'd0; 15271: data <= 'd0; 15272: data <= 'd0; 15273: data <= 'd0; 15274: data <= 'd0; 15275: data <= 'd2; 15276: data <= 'd4; 15277: data <= 'd7; 15278: data <= 'd2; 15279: data <= 'd0; 15280: data <= 'd0; 15281: data <= 'd0; 15282: data <= 'd0; 15283: data <= 'd2; 15284: data <= 'd4; 15285: data <= 'd4; 15286: data <= 'd2; 15287: data <= 'd0; 15288: data <= 'd0; 15289: data <= 'd0; 15290: data <= 'd0; 15291: data <= 'd0; 15292: data <= 'd0; 15293: data <= 'd0; 15294: data <= 'd0; 15295: data <= 'd0; 15296: data <= 'd0; 15297: data <= 'd0; 15298: data <= 'd0; 15299: data <= 'd0; 15300: data <= 'd0; 15301: data <= 'd0; 15302: data <= 'd0; 15303: data <= 'd0; 15304: data <= 'd0; 15305: data <= 'd0; 15306: data <= 'd0; 15307: data <= 'd2; 15308: data <= 'd2; 15309: data <= 'd2; 15310: data <= 'd0; 15311: data <= 'd0; 15312: data <= 'd0; 15313: data <= 'd0; 15314: data <= 'd0; 15315: data <= 'd0; 15316: data <= 'd2; 15317: data <= 'd2; 15318: data <= 'd2; 15319: data <= 'd0; 15320: data <= 'd0; 15321: data <= 'd0; 15322: data <= 'd0; 15323: data <= 'd0; 15324: data <= 'd0; 15325: data <= 'd0; 15326: data <= 'd0; 15327: data <= 'd0; 15328: data <= 'd0; 15329: data <= 'd0; 15330: data <= 'd0; 15331: data <= 'd0; 15332: data <= 'd0; 15333: data <= 'd0; 15334: data <= 'd0; 15335: data <= 'd0; 15336: data <= 'd0; 15337: data <= 'd0; 15338: data <= 'd0; 15339: data <= 'd0; 15340: data <= 'd0; 15341: data <= 'd0; 15342: data <= 'd0; 15343: data <= 'd0; 15344: data <= 'd0; 15345: data <= 'd0; 15346: data <= 'd0; 15347: data <= 'd0; 15348: data <= 'd0; 15349: data <= 'd0; 15350: data <= 'd0; 15351: data <= 'd0; 15352: data <= 'd0; 15353: data <= 'd0; 15354: data <= 'd0; 15355: data <= 'd0; 15356: data <= 'd0; 15357: data <= 'd0; 15358: data <= 'd0; 15359: data <= 'd0; 15360: data <= 'd0; 15361: data <= 'd0; 15362: data <= 'd0; 15363: data <= 'd0; 15364: data <= 'd0; 15365: data <= 'd0; 15366: data <= 'd0; 15367: data <= 'd0; 15368: data <= 'd0; 15369: data <= 'd0; 15370: data <= 'd0; 15371: data <= 'd0; 15372: data <= 'd0; 15373: data <= 'd0; 15374: data <= 'd0; 15375: data <= 'd0; 15376: data <= 'd0; 15377: data <= 'd0; 15378: data <= 'd0; 15379: data <= 'd0; 15380: data <= 'd0; 15381: data <= 'd0; 15382: data <= 'd0; 15383: data <= 'd0; 15384: data <= 'd0; 15385: data <= 'd0; 15386: data <= 'd0; 15387: data <= 'd0; 15388: data <= 'd0; 15389: data <= 'd0; 15390: data <= 'd0; 15391: data <= 'd0; 15392: data <= 'd0; 15393: data <= 'd0; 15394: data <= 'd0; 15395: data <= 'd0; 15396: data <= 'd0; 15397: data <= 'd0; 15398: data <= 'd0; 15399: data <= 'd0; 15400: data <= 'd0; 15401: data <= 'd0; 15402: data <= 'd0; 15403: data <= 'd0; 15404: data <= 'd0; 15405: data <= 'd0; 15406: data <= 'd0; 15407: data <= 'd0; 15408: data <= 'd0; 15409: data <= 'd0; 15410: data <= 'd0; 15411: data <= 'd0; 15412: data <= 'd0; 15413: data <= 'd0; 15414: data <= 'd0; 15415: data <= 'd0; 15416: data <= 'd0; 15417: data <= 'd0; 15418: data <= 'd0; 15419: data <= 'd0; 15420: data <= 'd0; 15421: data <= 'd0; 15422: data <= 'd0; 15423: data <= 'd0; 15424: data <= 'd0; 15425: data <= 'd0; 15426: data <= 'd0; 15427: data <= 'd0; 15428: data <= 'd0; 15429: data <= 'd0; 15430: data <= 'd0; 15431: data <= 'd0; 15432: data <= 'd0; 15433: data <= 'd0; 15434: data <= 'd0; 15435: data <= 'd0; 15436: data <= 'd0; 15437: data <= 'd0; 15438: data <= 'd0; 15439: data <= 'd0; 15440: data <= 'd0; 15441: data <= 'd0; 15442: data <= 'd0; 15443: data <= 'd0; 15444: data <= 'd0; 15445: data <= 'd0; 15446: data <= 'd0; 15447: data <= 'd0; 15448: data <= 'd0; 15449: data <= 'd0; 15450: data <= 'd0; 15451: data <= 'd0; 15452: data <= 'd0; 15453: data <= 'd0; 15454: data <= 'd0; 15455: data <= 'd0; 15456: data <= 'd0; 15457: data <= 'd0; 15458: data <= 'd0; 15459: data <= 'd0; 15460: data <= 'd0; 15461: data <= 'd0; 15462: data <= 'd0; 15463: data <= 'd0; 15464: data <= 'd0; 15465: data <= 'd0; 15466: data <= 'd0; 15467: data <= 'd0; 15468: data <= 'd0; 15469: data <= 'd0; 15470: data <= 'd0; 15471: data <= 'd0; 15472: data <= 'd0; 15473: data <= 'd0; 15474: data <= 'd0; 15475: data <= 'd0; 15476: data <= 'd0; 15477: data <= 'd0; 15478: data <= 'd0; 15479: data <= 'd0; 15480: data <= 'd0; 15481: data <= 'd0; 15482: data <= 'd0; 15483: data <= 'd0; 15484: data <= 'd0; 15485: data <= 'd0; 15486: data <= 'd0; 15487: data <= 'd0; 15488: data <= 'd0; 15489: data <= 'd0; 15490: data <= 'd0; 15491: data <= 'd0; 15492: data <= 'd0; 15493: data <= 'd0; 15494: data <= 'd0; 15495: data <= 'd0; 15496: data <= 'd0; 15497: data <= 'd0; 15498: data <= 'd0; 15499: data <= 'd0; 15500: data <= 'd0; 15501: data <= 'd0; 15502: data <= 'd0; 15503: data <= 'd0; 15504: data <= 'd0; 15505: data <= 'd0; 15506: data <= 'd0; 15507: data <= 'd0; 15508: data <= 'd0; 15509: data <= 'd0; 15510: data <= 'd0; 15511: data <= 'd0; 15512: data <= 'd0; 15513: data <= 'd0; 15514: data <= 'd0; 15515: data <= 'd0; 15516: data <= 'd0; 15517: data <= 'd0; 15518: data <= 'd0; 15519: data <= 'd0; 15520: data <= 'd0; 15521: data <= 'd0; 15522: data <= 'd0; 15523: data <= 'd0; 15524: data <= 'd0; 15525: data <= 'd0; 15526: data <= 'd0; 15527: data <= 'd0; 15528: data <= 'd0; 15529: data <= 'd0; 15530: data <= 'd0; 15531: data <= 'd0; 15532: data <= 'd0; 15533: data <= 'd0; 15534: data <= 'd0; 15535: data <= 'd0; 15536: data <= 'd0; 15537: data <= 'd0; 15538: data <= 'd0; 15539: data <= 'd0; 15540: data <= 'd0; 15541: data <= 'd0; 15542: data <= 'd0; 15543: data <= 'd0; 15544: data <= 'd0; 15545: data <= 'd0; 15546: data <= 'd0; 15547: data <= 'd0; 15548: data <= 'd0; 15549: data <= 'd0; 15550: data <= 'd0; 15551: data <= 'd0; 15552: data <= 'd0; 15553: data <= 'd0; 15554: data <= 'd0; 15555: data <= 'd0; 15556: data <= 'd0; 15557: data <= 'd0; 15558: data <= 'd0; 15559: data <= 'd0; 15560: data <= 'd0; 15561: data <= 'd0; 15562: data <= 'd0; 15563: data <= 'd0; 15564: data <= 'd0; 15565: data <= 'd0; 15566: data <= 'd0; 15567: data <= 'd0; 15568: data <= 'd0; 15569: data <= 'd0; 15570: data <= 'd0; 15571: data <= 'd0; 15572: data <= 'd0; 15573: data <= 'd0; 15574: data <= 'd0; 15575: data <= 'd0; 15576: data <= 'd0; 15577: data <= 'd0; 15578: data <= 'd0; 15579: data <= 'd0; 15580: data <= 'd0; 15581: data <= 'd0; 15582: data <= 'd0; 15583: data <= 'd0; 15584: data <= 'd0; 15585: data <= 'd0; 15586: data <= 'd0; 15587: data <= 'd0; 15588: data <= 'd0; 15589: data <= 'd0; 15590: data <= 'd0; 15591: data <= 'd0; 15592: data <= 'd0; 15593: data <= 'd0; 15594: data <= 'd0; 15595: data <= 'd0; 15596: data <= 'd0; 15597: data <= 'd0; 15598: data <= 'd0; 15599: data <= 'd0; 15600: data <= 'd0; 15601: data <= 'd0; 15602: data <= 'd0; 15603: data <= 'd0; 15604: data <= 'd0; 15605: data <= 'd0; 15606: data <= 'd0; 15607: data <= 'd0; 15608: data <= 'd0; 15609: data <= 'd0; 15610: data <= 'd0; 15611: data <= 'd0; 15612: data <= 'd0; 15613: data <= 'd0; 15614: data <= 'd0; 15615: data <= 'd0; 15616: data <= 'd0; 15617: data <= 'd0; 15618: data <= 'd0; 15619: data <= 'd0; 15620: data <= 'd0; 15621: data <= 'd0; 15622: data <= 'd0; 15623: data <= 'd0; 15624: data <= 'd0; 15625: data <= 'd0; 15626: data <= 'd0; 15627: data <= 'd0; 15628: data <= 'd0; 15629: data <= 'd0; 15630: data <= 'd0; 15631: data <= 'd0; 15632: data <= 'd0; 15633: data <= 'd0; 15634: data <= 'd0; 15635: data <= 'd0; 15636: data <= 'd0; 15637: data <= 'd0; 15638: data <= 'd0; 15639: data <= 'd0; 15640: data <= 'd0; 15641: data <= 'd0; 15642: data <= 'd0; 15643: data <= 'd0; 15644: data <= 'd0; 15645: data <= 'd0; 15646: data <= 'd0; 15647: data <= 'd0; 15648: data <= 'd0; 15649: data <= 'd0; 15650: data <= 'd0; 15651: data <= 'd0; 15652: data <= 'd0; 15653: data <= 'd0; 15654: data <= 'd0; 15655: data <= 'd0; 15656: data <= 'd0; 15657: data <= 'd0; 15658: data <= 'd0; 15659: data <= 'd0; 15660: data <= 'd0; 15661: data <= 'd2; 15662: data <= 'd2; 15663: data <= 'd2; 15664: data <= 'd2; 15665: data <= 'd2; 15666: data <= 'd2; 15667: data <= 'd0; 15668: data <= 'd0; 15669: data <= 'd0; 15670: data <= 'd0; 15671: data <= 'd0; 15672: data <= 'd0; 15673: data <= 'd0; 15674: data <= 'd0; 15675: data <= 'd0; 15676: data <= 'd0; 15677: data <= 'd0; 15678: data <= 'd0; 15679: data <= 'd0; 15680: data <= 'd0; 15681: data <= 'd0; 15682: data <= 'd0; 15683: data <= 'd0; 15684: data <= 'd0; 15685: data <= 'd0; 15686: data <= 'd0; 15687: data <= 'd0; 15688: data <= 'd0; 15689: data <= 'd0; 15690: data <= 'd0; 15691: data <= 'd2; 15692: data <= 'd2; 15693: data <= 'd6; 15694: data <= 'd6; 15695: data <= 'd6; 15696: data <= 'd6; 15697: data <= 'd6; 15698: data <= 'd6; 15699: data <= 'd2; 15700: data <= 'd2; 15701: data <= 'd0; 15702: data <= 'd0; 15703: data <= 'd0; 15704: data <= 'd0; 15705: data <= 'd0; 15706: data <= 'd0; 15707: data <= 'd0; 15708: data <= 'd0; 15709: data <= 'd0; 15710: data <= 'd0; 15711: data <= 'd0; 15712: data <= 'd0; 15713: data <= 'd0; 15714: data <= 'd0; 15715: data <= 'd0; 15716: data <= 'd0; 15717: data <= 'd0; 15718: data <= 'd0; 15719: data <= 'd0; 15720: data <= 'd0; 15721: data <= 'd0; 15722: data <= 'd2; 15723: data <= 'd1; 15724: data <= 'd3; 15725: data <= 'd6; 15726: data <= 'd6; 15727: data <= 'd6; 15728: data <= 'd6; 15729: data <= 'd6; 15730: data <= 'd6; 15731: data <= 'd6; 15732: data <= 'd3; 15733: data <= 'd2; 15734: data <= 'd0; 15735: data <= 'd0; 15736: data <= 'd0; 15737: data <= 'd0; 15738: data <= 'd0; 15739: data <= 'd0; 15740: data <= 'd0; 15741: data <= 'd0; 15742: data <= 'd0; 15743: data <= 'd0; 15744: data <= 'd0; 15745: data <= 'd0; 15746: data <= 'd0; 15747: data <= 'd0; 15748: data <= 'd0; 15749: data <= 'd0; 15750: data <= 'd0; 15751: data <= 'd0; 15752: data <= 'd0; 15753: data <= 'd2; 15754: data <= 'd1; 15755: data <= 'd1; 15756: data <= 'd1; 15757: data <= 'd3; 15758: data <= 'd6; 15759: data <= 'd6; 15760: data <= 'd6; 15761: data <= 'd6; 15762: data <= 'd6; 15763: data <= 'd3; 15764: data <= 'd1; 15765: data <= 'd1; 15766: data <= 'd2; 15767: data <= 'd0; 15768: data <= 'd0; 15769: data <= 'd0; 15770: data <= 'd0; 15771: data <= 'd0; 15772: data <= 'd0; 15773: data <= 'd0; 15774: data <= 'd0; 15775: data <= 'd0; 15776: data <= 'd0; 15777: data <= 'd0; 15778: data <= 'd0; 15779: data <= 'd0; 15780: data <= 'd0; 15781: data <= 'd0; 15782: data <= 'd0; 15783: data <= 'd0; 15784: data <= 'd0; 15785: data <= 'd2; 15786: data <= 'd1; 15787: data <= 'd1; 15788: data <= 'd5; 15789: data <= 'd5; 15790: data <= 'd5; 15791: data <= 'd1; 15792: data <= 'd1; 15793: data <= 'd1; 15794: data <= 'd1; 15795: data <= 'd1; 15796: data <= 'd5; 15797: data <= 'd5; 15798: data <= 'd2; 15799: data <= 'd0; 15800: data <= 'd0; 15801: data <= 'd0; 15802: data <= 'd0; 15803: data <= 'd0; 15804: data <= 'd0; 15805: data <= 'd0; 15806: data <= 'd0; 15807: data <= 'd0; 15808: data <= 'd0; 15809: data <= 'd0; 15810: data <= 'd0; 15811: data <= 'd0; 15812: data <= 'd0; 15813: data <= 'd0; 15814: data <= 'd0; 15815: data <= 'd0; 15816: data <= 'd2; 15817: data <= 'd1; 15818: data <= 'd5; 15819: data <= 'd5; 15820: data <= 'd3; 15821: data <= 'd6; 15822: data <= 'd6; 15823: data <= 'd6; 15824: data <= 'd6; 15825: data <= 'd6; 15826: data <= 'd6; 15827: data <= 'd6; 15828: data <= 'd6; 15829: data <= 'd3; 15830: data <= 'd5; 15831: data <= 'd2; 15832: data <= 'd0; 15833: data <= 'd0; 15834: data <= 'd0; 15835: data <= 'd0; 15836: data <= 'd0; 15837: data <= 'd0; 15838: data <= 'd0; 15839: data <= 'd0; 15840: data <= 'd0; 15841: data <= 'd0; 15842: data <= 'd0; 15843: data <= 'd0; 15844: data <= 'd0; 15845: data <= 'd0; 15846: data <= 'd0; 15847: data <= 'd0; 15848: data <= 'd2; 15849: data <= 'd5; 15850: data <= 'd3; 15851: data <= 'd6; 15852: data <= 'd3; 15853: data <= 'd1; 15854: data <= 'd1; 15855: data <= 'd1; 15856: data <= 'd1; 15857: data <= 'd1; 15858: data <= 'd1; 15859: data <= 'd1; 15860: data <= 'd1; 15861: data <= 'd1; 15862: data <= 'd3; 15863: data <= 'd2; 15864: data <= 'd0; 15865: data <= 'd0; 15866: data <= 'd0; 15867: data <= 'd0; 15868: data <= 'd0; 15869: data <= 'd0; 15870: data <= 'd0; 15871: data <= 'd0; 15872: data <= 'd0; 15873: data <= 'd0; 15874: data <= 'd0; 15875: data <= 'd0; 15876: data <= 'd0; 15877: data <= 'd0; 15878: data <= 'd0; 15879: data <= 'd0; 15880: data <= 'd2; 15881: data <= 'd5; 15882: data <= 'd3; 15883: data <= 'd1; 15884: data <= 'd1; 15885: data <= 'd1; 15886: data <= 'd5; 15887: data <= 'd5; 15888: data <= 'd5; 15889: data <= 'd5; 15890: data <= 'd5; 15891: data <= 'd5; 15892: data <= 'd5; 15893: data <= 'd1; 15894: data <= 'd1; 15895: data <= 'd2; 15896: data <= 'd0; 15897: data <= 'd0; 15898: data <= 'd0; 15899: data <= 'd0; 15900: data <= 'd0; 15901: data <= 'd0; 15902: data <= 'd0; 15903: data <= 'd0; 15904: data <= 'd0; 15905: data <= 'd0; 15906: data <= 'd0; 15907: data <= 'd0; 15908: data <= 'd0; 15909: data <= 'd0; 15910: data <= 'd0; 15911: data <= 'd0; 15912: data <= 'd2; 15913: data <= 'd6; 15914: data <= 'd1; 15915: data <= 'd5; 15916: data <= 'd2; 15917: data <= 'd2; 15918: data <= 'd2; 15919: data <= 'd2; 15920: data <= 'd2; 15921: data <= 'd2; 15922: data <= 'd2; 15923: data <= 'd2; 15924: data <= 'd2; 15925: data <= 'd2; 15926: data <= 'd5; 15927: data <= 'd2; 15928: data <= 'd0; 15929: data <= 'd0; 15930: data <= 'd0; 15931: data <= 'd0; 15932: data <= 'd0; 15933: data <= 'd0; 15934: data <= 'd0; 15935: data <= 'd0; 15936: data <= 'd0; 15937: data <= 'd0; 15938: data <= 'd0; 15939: data <= 'd0; 15940: data <= 'd0; 15941: data <= 'd0; 15942: data <= 'd2; 15943: data <= 'd2; 15944: data <= 'd5; 15945: data <= 'd6; 15946: data <= 'd5; 15947: data <= 'd2; 15948: data <= 'd8; 15949: data <= 'd8; 15950: data <= 'd8; 15951: data <= 'd8; 15952: data <= 'd8; 15953: data <= 'd9; 15954: data <= 'd9; 15955: data <= 'd8; 15956: data <= 'd8; 15957: data <= 'd8; 15958: data <= 'd2; 15959: data <= 'd2; 15960: data <= 'd0; 15961: data <= 'd0; 15962: data <= 'd0; 15963: data <= 'd0; 15964: data <= 'd0; 15965: data <= 'd0; 15966: data <= 'd0; 15967: data <= 'd0; 15968: data <= 'd0; 15969: data <= 'd0; 15970: data <= 'd0; 15971: data <= 'd0; 15972: data <= 'd0; 15973: data <= 'd0; 15974: data <= 'd2; 15975: data <= 'd3; 15976: data <= 'd6; 15977: data <= 'd3; 15978: data <= 'd2; 15979: data <= 'd8; 15980: data <= 'd8; 15981: data <= 'd9; 15982: data <= 'd9; 15983: data <= 'd10; 15984: data <= 'd2; 15985: data <= 'd9; 15986: data <= 'd11; 15987: data <= 'd10; 15988: data <= 'd2; 15989: data <= 'd9; 15990: data <= 'd2; 15991: data <= 'd2; 15992: data <= 'd0; 15993: data <= 'd0; 15994: data <= 'd0; 15995: data <= 'd0; 15996: data <= 'd0; 15997: data <= 'd0; 15998: data <= 'd0; 15999: data <= 'd0; 16000: data <= 'd0; 16001: data <= 'd0; 16002: data <= 'd0; 16003: data <= 'd0; 16004: data <= 'd0; 16005: data <= 'd0; 16006: data <= 'd2; 16007: data <= 'd1; 16008: data <= 'd3; 16009: data <= 'd1; 16010: data <= 'd2; 16011: data <= 'd10; 16012: data <= 'd10; 16013: data <= 'd9; 16014: data <= 'd10; 16015: data <= 'd10; 16016: data <= 'd11; 16017: data <= 'd10; 16018: data <= 'd11; 16019: data <= 'd11; 16020: data <= 'd10; 16021: data <= 'd10; 16022: data <= 'd2; 16023: data <= 'd0; 16024: data <= 'd0; 16025: data <= 'd0; 16026: data <= 'd0; 16027: data <= 'd0; 16028: data <= 'd0; 16029: data <= 'd0; 16030: data <= 'd0; 16031: data <= 'd0; 16032: data <= 'd0; 16033: data <= 'd0; 16034: data <= 'd0; 16035: data <= 'd0; 16036: data <= 'd0; 16037: data <= 'd0; 16038: data <= 'd0; 16039: data <= 'd2; 16040: data <= 'd1; 16041: data <= 'd5; 16042: data <= 'd2; 16043: data <= 'd8; 16044: data <= 'd9; 16045: data <= 'd9; 16046: data <= 'd10; 16047: data <= 'd10; 16048: data <= 'd10; 16049: data <= 'd10; 16050: data <= 'd8; 16051: data <= 'd8; 16052: data <= 'd10; 16053: data <= 'd9; 16054: data <= 'd2; 16055: data <= 'd0; 16056: data <= 'd0; 16057: data <= 'd0; 16058: data <= 'd0; 16059: data <= 'd0; 16060: data <= 'd0; 16061: data <= 'd0; 16062: data <= 'd0; 16063: data <= 'd0; 16064: data <= 'd0; 16065: data <= 'd0; 16066: data <= 'd0; 16067: data <= 'd0; 16068: data <= 'd0; 16069: data <= 'd0; 16070: data <= 'd0; 16071: data <= 'd0; 16072: data <= 'd2; 16073: data <= 'd2; 16074: data <= 'd2; 16075: data <= 'd8; 16076: data <= 'd8; 16077: data <= 'd9; 16078: data <= 'd9; 16079: data <= 'd10; 16080: data <= 'd10; 16081: data <= 'd10; 16082: data <= 'd9; 16083: data <= 'd9; 16084: data <= 'd10; 16085: data <= 'd9; 16086: data <= 'd2; 16087: data <= 'd0; 16088: data <= 'd0; 16089: data <= 'd0; 16090: data <= 'd0; 16091: data <= 'd0; 16092: data <= 'd0; 16093: data <= 'd0; 16094: data <= 'd0; 16095: data <= 'd0; 16096: data <= 'd0; 16097: data <= 'd0; 16098: data <= 'd0; 16099: data <= 'd0; 16100: data <= 'd0; 16101: data <= 'd0; 16102: data <= 'd0; 16103: data <= 'd0; 16104: data <= 'd0; 16105: data <= 'd0; 16106: data <= 'd0; 16107: data <= 'd2; 16108: data <= 'd5; 16109: data <= 'd5; 16110: data <= 'd8; 16111: data <= 'd9; 16112: data <= 'd9; 16113: data <= 'd9; 16114: data <= 'd9; 16115: data <= 'd9; 16116: data <= 'd9; 16117: data <= 'd2; 16118: data <= 'd0; 16119: data <= 'd0; 16120: data <= 'd0; 16121: data <= 'd0; 16122: data <= 'd0; 16123: data <= 'd0; 16124: data <= 'd0; 16125: data <= 'd0; 16126: data <= 'd0; 16127: data <= 'd0; 16128: data <= 'd0; 16129: data <= 'd0; 16130: data <= 'd0; 16131: data <= 'd0; 16132: data <= 'd0; 16133: data <= 'd0; 16134: data <= 'd0; 16135: data <= 'd0; 16136: data <= 'd0; 16137: data <= 'd0; 16138: data <= 'd2; 16139: data <= 'd7; 16140: data <= 'd1; 16141: data <= 'd1; 16142: data <= 'd1; 16143: data <= 'd3; 16144: data <= 'd3; 16145: data <= 'd3; 16146: data <= 'd5; 16147: data <= 'd5; 16148: data <= 'd3; 16149: data <= 'd1; 16150: data <= 'd2; 16151: data <= 'd0; 16152: data <= 'd0; 16153: data <= 'd0; 16154: data <= 'd0; 16155: data <= 'd0; 16156: data <= 'd0; 16157: data <= 'd0; 16158: data <= 'd0; 16159: data <= 'd0; 16160: data <= 'd0; 16161: data <= 'd0; 16162: data <= 'd0; 16163: data <= 'd0; 16164: data <= 'd0; 16165: data <= 'd0; 16166: data <= 'd0; 16167: data <= 'd0; 16168: data <= 'd0; 16169: data <= 'd0; 16170: data <= 'd2; 16171: data <= 'd7; 16172: data <= 'd7; 16173: data <= 'd1; 16174: data <= 'd1; 16175: data <= 'd3; 16176: data <= 'd3; 16177: data <= 'd3; 16178: data <= 'd1; 16179: data <= 'd1; 16180: data <= 'd3; 16181: data <= 'd1; 16182: data <= 'd2; 16183: data <= 'd0; 16184: data <= 'd0; 16185: data <= 'd0; 16186: data <= 'd0; 16187: data <= 'd0; 16188: data <= 'd0; 16189: data <= 'd0; 16190: data <= 'd0; 16191: data <= 'd0; 16192: data <= 'd0; 16193: data <= 'd0; 16194: data <= 'd0; 16195: data <= 'd0; 16196: data <= 'd0; 16197: data <= 'd0; 16198: data <= 'd0; 16199: data <= 'd0; 16200: data <= 'd0; 16201: data <= 'd2; 16202: data <= 'd9; 16203: data <= 'd9; 16204: data <= 'd7; 16205: data <= 'd1; 16206: data <= 'd1; 16207: data <= 'd1; 16208: data <= 'd3; 16209: data <= 'd3; 16210: data <= 'd1; 16211: data <= 'd1; 16212: data <= 'd1; 16213: data <= 'd1; 16214: data <= 'd8; 16215: data <= 'd2; 16216: data <= 'd0; 16217: data <= 'd0; 16218: data <= 'd0; 16219: data <= 'd0; 16220: data <= 'd0; 16221: data <= 'd0; 16222: data <= 'd0; 16223: data <= 'd0; 16224: data <= 'd0; 16225: data <= 'd0; 16226: data <= 'd0; 16227: data <= 'd0; 16228: data <= 'd0; 16229: data <= 'd0; 16230: data <= 'd0; 16231: data <= 'd0; 16232: data <= 'd0; 16233: data <= 'd2; 16234: data <= 'd9; 16235: data <= 'd9; 16236: data <= 'd2; 16237: data <= 'd2; 16238: data <= 'd2; 16239: data <= 'd2; 16240: data <= 'd2; 16241: data <= 'd5; 16242: data <= 'd5; 16243: data <= 'd5; 16244: data <= 'd2; 16245: data <= 'd2; 16246: data <= 'd8; 16247: data <= 'd2; 16248: data <= 'd0; 16249: data <= 'd0; 16250: data <= 'd0; 16251: data <= 'd0; 16252: data <= 'd0; 16253: data <= 'd0; 16254: data <= 'd0; 16255: data <= 'd0; 16256: data <= 'd0; 16257: data <= 'd0; 16258: data <= 'd0; 16259: data <= 'd0; 16260: data <= 'd0; 16261: data <= 'd0; 16262: data <= 'd0; 16263: data <= 'd0; 16264: data <= 'd0; 16265: data <= 'd0; 16266: data <= 'd2; 16267: data <= 'd2; 16268: data <= 'd2; 16269: data <= 'd1; 16270: data <= 'd1; 16271: data <= 'd3; 16272: data <= 'd5; 16273: data <= 'd1; 16274: data <= 'd3; 16275: data <= 'd3; 16276: data <= 'd3; 16277: data <= 'd2; 16278: data <= 'd2; 16279: data <= 'd0; 16280: data <= 'd0; 16281: data <= 'd0; 16282: data <= 'd0; 16283: data <= 'd0; 16284: data <= 'd0; 16285: data <= 'd0; 16286: data <= 'd0; 16287: data <= 'd0; 16288: data <= 'd0; 16289: data <= 'd0; 16290: data <= 'd0; 16291: data <= 'd0; 16292: data <= 'd0; 16293: data <= 'd0; 16294: data <= 'd0; 16295: data <= 'd0; 16296: data <= 'd0; 16297: data <= 'd0; 16298: data <= 'd0; 16299: data <= 'd0; 16300: data <= 'd0; 16301: data <= 'd2; 16302: data <= 'd4; 16303: data <= 'd7; 16304: data <= 'd2; 16305: data <= 'd2; 16306: data <= 'd5; 16307: data <= 'd5; 16308: data <= 'd4; 16309: data <= 'd2; 16310: data <= 'd0; 16311: data <= 'd0; 16312: data <= 'd0; 16313: data <= 'd0; 16314: data <= 'd0; 16315: data <= 'd0; 16316: data <= 'd0; 16317: data <= 'd0; 16318: data <= 'd0; 16319: data <= 'd0; 16320: data <= 'd0; 16321: data <= 'd0; 16322: data <= 'd0; 16323: data <= 'd0; 16324: data <= 'd0; 16325: data <= 'd0; 16326: data <= 'd0; 16327: data <= 'd0; 16328: data <= 'd0; 16329: data <= 'd0; 16330: data <= 'd0; 16331: data <= 'd0; 16332: data <= 'd0; 16333: data <= 'd2; 16334: data <= 'd2; 16335: data <= 'd2; 16336: data <= 'd0; 16337: data <= 'd2; 16338: data <= 'd4; 16339: data <= 'd4; 16340: data <= 'd2; 16341: data <= 'd0; 16342: data <= 'd0; 16343: data <= 'd0; 16344: data <= 'd0; 16345: data <= 'd0; 16346: data <= 'd0; 16347: data <= 'd0; 16348: data <= 'd0; 16349: data <= 'd0; 16350: data <= 'd0; 16351: data <= 'd0; 16352: data <= 'd0; 16353: data <= 'd0; 16354: data <= 'd0; 16355: data <= 'd0; 16356: data <= 'd0; 16357: data <= 'd0; 16358: data <= 'd0; 16359: data <= 'd0; 16360: data <= 'd0; 16361: data <= 'd0; 16362: data <= 'd0; 16363: data <= 'd0; 16364: data <= 'd0; 16365: data <= 'd0; 16366: data <= 'd0; 16367: data <= 'd0; 16368: data <= 'd0; 16369: data <= 'd2; 16370: data <= 'd2; 16371: data <= 'd2; 16372: data <= 'd0; 16373: data <= 'd0; 16374: data <= 'd0; 16375: data <= 'd0; 16376: data <= 'd0; 16377: data <= 'd0; 16378: data <= 'd0; 16379: data <= 'd0; 16380: data <= 'd0; 16381: data <= 'd0; 16382: data <= 'd0; 16383: data <= 'd0; 16384: data <= 'd0; 16385: data <= 'd0; 16386: data <= 'd0; 16387: data <= 'd0; 16388: data <= 'd0; 16389: data <= 'd0; 16390: data <= 'd0; 16391: data <= 'd0; 16392: data <= 'd0; 16393: data <= 'd0; 16394: data <= 'd0; 16395: data <= 'd0; 16396: data <= 'd0; 16397: data <= 'd0; 16398: data <= 'd0; 16399: data <= 'd0; 16400: data <= 'd0; 16401: data <= 'd0; 16402: data <= 'd0; 16403: data <= 'd0; 16404: data <= 'd0; 16405: data <= 'd0; 16406: data <= 'd0; 16407: data <= 'd0; 16408: data <= 'd0; 16409: data <= 'd0; 16410: data <= 'd0; 16411: data <= 'd0; 16412: data <= 'd0; 16413: data <= 'd0; 16414: data <= 'd0; 16415: data <= 'd0; 16416: data <= 'd0; 16417: data <= 'd0; 16418: data <= 'd0; 16419: data <= 'd0; 16420: data <= 'd0; 16421: data <= 'd0; 16422: data <= 'd0; 16423: data <= 'd0; 16424: data <= 'd0; 16425: data <= 'd0; 16426: data <= 'd0; 16427: data <= 'd0; 16428: data <= 'd0; 16429: data <= 'd0; 16430: data <= 'd0; 16431: data <= 'd0; 16432: data <= 'd0; 16433: data <= 'd0; 16434: data <= 'd0; 16435: data <= 'd0; 16436: data <= 'd0; 16437: data <= 'd0; 16438: data <= 'd0; 16439: data <= 'd0; 16440: data <= 'd0; 16441: data <= 'd0; 16442: data <= 'd0; 16443: data <= 'd0; 16444: data <= 'd0; 16445: data <= 'd0; 16446: data <= 'd0; 16447: data <= 'd0; 16448: data <= 'd0; 16449: data <= 'd0; 16450: data <= 'd0; 16451: data <= 'd0; 16452: data <= 'd0; 16453: data <= 'd0; 16454: data <= 'd0; 16455: data <= 'd0; 16456: data <= 'd0; 16457: data <= 'd0; 16458: data <= 'd0; 16459: data <= 'd0; 16460: data <= 'd0; 16461: data <= 'd0; 16462: data <= 'd0; 16463: data <= 'd0; 16464: data <= 'd0; 16465: data <= 'd0; 16466: data <= 'd0; 16467: data <= 'd0; 16468: data <= 'd0; 16469: data <= 'd0; 16470: data <= 'd0; 16471: data <= 'd0; 16472: data <= 'd0; 16473: data <= 'd0; 16474: data <= 'd0; 16475: data <= 'd0; 16476: data <= 'd0; 16477: data <= 'd0; 16478: data <= 'd0; 16479: data <= 'd0; 16480: data <= 'd0; 16481: data <= 'd0; 16482: data <= 'd0; 16483: data <= 'd0; 16484: data <= 'd0; 16485: data <= 'd0; 16486: data <= 'd0; 16487: data <= 'd0; 16488: data <= 'd0; 16489: data <= 'd0; 16490: data <= 'd0; 16491: data <= 'd0; 16492: data <= 'd0; 16493: data <= 'd0; 16494: data <= 'd0; 16495: data <= 'd0; 16496: data <= 'd0; 16497: data <= 'd0; 16498: data <= 'd0; 16499: data <= 'd0; 16500: data <= 'd0; 16501: data <= 'd0; 16502: data <= 'd0; 16503: data <= 'd0; 16504: data <= 'd0; 16505: data <= 'd0; 16506: data <= 'd0; 16507: data <= 'd0; 16508: data <= 'd0; 16509: data <= 'd0; 16510: data <= 'd0; 16511: data <= 'd0; 16512: data <= 'd0; 16513: data <= 'd0; 16514: data <= 'd0; 16515: data <= 'd0; 16516: data <= 'd0; 16517: data <= 'd0; 16518: data <= 'd0; 16519: data <= 'd0; 16520: data <= 'd0; 16521: data <= 'd0; 16522: data <= 'd0; 16523: data <= 'd0; 16524: data <= 'd0; 16525: data <= 'd0; 16526: data <= 'd0; 16527: data <= 'd0; 16528: data <= 'd0; 16529: data <= 'd0; 16530: data <= 'd0; 16531: data <= 'd0; 16532: data <= 'd0; 16533: data <= 'd0; 16534: data <= 'd0; 16535: data <= 'd0; 16536: data <= 'd0; 16537: data <= 'd0; 16538: data <= 'd0; 16539: data <= 'd0; 16540: data <= 'd0; 16541: data <= 'd0; 16542: data <= 'd0; 16543: data <= 'd0; 16544: data <= 'd0; 16545: data <= 'd0; 16546: data <= 'd0; 16547: data <= 'd0; 16548: data <= 'd0; 16549: data <= 'd0; 16550: data <= 'd0; 16551: data <= 'd0; 16552: data <= 'd0; 16553: data <= 'd0; 16554: data <= 'd0; 16555: data <= 'd0; 16556: data <= 'd0; 16557: data <= 'd0; 16558: data <= 'd0; 16559: data <= 'd0; 16560: data <= 'd0; 16561: data <= 'd0; 16562: data <= 'd0; 16563: data <= 'd0; 16564: data <= 'd0; 16565: data <= 'd0; 16566: data <= 'd0; 16567: data <= 'd0; 16568: data <= 'd0; 16569: data <= 'd0; 16570: data <= 'd0; 16571: data <= 'd0; 16572: data <= 'd0; 16573: data <= 'd0; 16574: data <= 'd0; 16575: data <= 'd0; 16576: data <= 'd0; 16577: data <= 'd0; 16578: data <= 'd0; 16579: data <= 'd0; 16580: data <= 'd0; 16581: data <= 'd0; 16582: data <= 'd0; 16583: data <= 'd0; 16584: data <= 'd0; 16585: data <= 'd0; 16586: data <= 'd0; 16587: data <= 'd0; 16588: data <= 'd0; 16589: data <= 'd0; 16590: data <= 'd0; 16591: data <= 'd0; 16592: data <= 'd0; 16593: data <= 'd0; 16594: data <= 'd0; 16595: data <= 'd0; 16596: data <= 'd0; 16597: data <= 'd0; 16598: data <= 'd0; 16599: data <= 'd0; 16600: data <= 'd0; 16601: data <= 'd0; 16602: data <= 'd0; 16603: data <= 'd0; 16604: data <= 'd0; 16605: data <= 'd0; 16606: data <= 'd0; 16607: data <= 'd0; 16608: data <= 'd0; 16609: data <= 'd0; 16610: data <= 'd0; 16611: data <= 'd0; 16612: data <= 'd0; 16613: data <= 'd0; 16614: data <= 'd0; 16615: data <= 'd0; 16616: data <= 'd0; 16617: data <= 'd0; 16618: data <= 'd0; 16619: data <= 'd0; 16620: data <= 'd0; 16621: data <= 'd0; 16622: data <= 'd0; 16623: data <= 'd0; 16624: data <= 'd0; 16625: data <= 'd0; 16626: data <= 'd0; 16627: data <= 'd0; 16628: data <= 'd0; 16629: data <= 'd0; 16630: data <= 'd0; 16631: data <= 'd0; 16632: data <= 'd0; 16633: data <= 'd0; 16634: data <= 'd0; 16635: data <= 'd0; 16636: data <= 'd0; 16637: data <= 'd0; 16638: data <= 'd0; 16639: data <= 'd0; 16640: data <= 'd0; 16641: data <= 'd0; 16642: data <= 'd0; 16643: data <= 'd0; 16644: data <= 'd0; 16645: data <= 'd0; 16646: data <= 'd0; 16647: data <= 'd0; 16648: data <= 'd0; 16649: data <= 'd0; 16650: data <= 'd0; 16651: data <= 'd0; 16652: data <= 'd0; 16653: data <= 'd2; 16654: data <= 'd2; 16655: data <= 'd2; 16656: data <= 'd2; 16657: data <= 'd2; 16658: data <= 'd2; 16659: data <= 'd0; 16660: data <= 'd0; 16661: data <= 'd0; 16662: data <= 'd0; 16663: data <= 'd0; 16664: data <= 'd0; 16665: data <= 'd0; 16666: data <= 'd0; 16667: data <= 'd0; 16668: data <= 'd0; 16669: data <= 'd0; 16670: data <= 'd0; 16671: data <= 'd0; 16672: data <= 'd0; 16673: data <= 'd0; 16674: data <= 'd0; 16675: data <= 'd0; 16676: data <= 'd0; 16677: data <= 'd0; 16678: data <= 'd0; 16679: data <= 'd0; 16680: data <= 'd0; 16681: data <= 'd0; 16682: data <= 'd0; 16683: data <= 'd2; 16684: data <= 'd2; 16685: data <= 'd6; 16686: data <= 'd6; 16687: data <= 'd6; 16688: data <= 'd6; 16689: data <= 'd6; 16690: data <= 'd6; 16691: data <= 'd2; 16692: data <= 'd2; 16693: data <= 'd0; 16694: data <= 'd0; 16695: data <= 'd0; 16696: data <= 'd0; 16697: data <= 'd0; 16698: data <= 'd0; 16699: data <= 'd0; 16700: data <= 'd0; 16701: data <= 'd0; 16702: data <= 'd0; 16703: data <= 'd0; 16704: data <= 'd0; 16705: data <= 'd0; 16706: data <= 'd0; 16707: data <= 'd0; 16708: data <= 'd0; 16709: data <= 'd0; 16710: data <= 'd0; 16711: data <= 'd0; 16712: data <= 'd0; 16713: data <= 'd0; 16714: data <= 'd2; 16715: data <= 'd1; 16716: data <= 'd3; 16717: data <= 'd6; 16718: data <= 'd6; 16719: data <= 'd6; 16720: data <= 'd6; 16721: data <= 'd6; 16722: data <= 'd6; 16723: data <= 'd6; 16724: data <= 'd3; 16725: data <= 'd2; 16726: data <= 'd0; 16727: data <= 'd0; 16728: data <= 'd0; 16729: data <= 'd0; 16730: data <= 'd0; 16731: data <= 'd0; 16732: data <= 'd0; 16733: data <= 'd0; 16734: data <= 'd0; 16735: data <= 'd0; 16736: data <= 'd0; 16737: data <= 'd0; 16738: data <= 'd0; 16739: data <= 'd0; 16740: data <= 'd0; 16741: data <= 'd0; 16742: data <= 'd0; 16743: data <= 'd0; 16744: data <= 'd0; 16745: data <= 'd2; 16746: data <= 'd1; 16747: data <= 'd1; 16748: data <= 'd1; 16749: data <= 'd3; 16750: data <= 'd6; 16751: data <= 'd6; 16752: data <= 'd6; 16753: data <= 'd6; 16754: data <= 'd6; 16755: data <= 'd3; 16756: data <= 'd1; 16757: data <= 'd1; 16758: data <= 'd2; 16759: data <= 'd0; 16760: data <= 'd0; 16761: data <= 'd0; 16762: data <= 'd0; 16763: data <= 'd0; 16764: data <= 'd0; 16765: data <= 'd0; 16766: data <= 'd0; 16767: data <= 'd0; 16768: data <= 'd0; 16769: data <= 'd0; 16770: data <= 'd0; 16771: data <= 'd0; 16772: data <= 'd0; 16773: data <= 'd0; 16774: data <= 'd0; 16775: data <= 'd0; 16776: data <= 'd0; 16777: data <= 'd2; 16778: data <= 'd1; 16779: data <= 'd1; 16780: data <= 'd5; 16781: data <= 'd5; 16782: data <= 'd5; 16783: data <= 'd1; 16784: data <= 'd1; 16785: data <= 'd1; 16786: data <= 'd1; 16787: data <= 'd1; 16788: data <= 'd5; 16789: data <= 'd5; 16790: data <= 'd2; 16791: data <= 'd0; 16792: data <= 'd0; 16793: data <= 'd0; 16794: data <= 'd0; 16795: data <= 'd0; 16796: data <= 'd0; 16797: data <= 'd0; 16798: data <= 'd0; 16799: data <= 'd0; 16800: data <= 'd0; 16801: data <= 'd0; 16802: data <= 'd0; 16803: data <= 'd0; 16804: data <= 'd0; 16805: data <= 'd0; 16806: data <= 'd0; 16807: data <= 'd0; 16808: data <= 'd2; 16809: data <= 'd1; 16810: data <= 'd5; 16811: data <= 'd5; 16812: data <= 'd3; 16813: data <= 'd6; 16814: data <= 'd6; 16815: data <= 'd6; 16816: data <= 'd6; 16817: data <= 'd6; 16818: data <= 'd6; 16819: data <= 'd6; 16820: data <= 'd6; 16821: data <= 'd3; 16822: data <= 'd5; 16823: data <= 'd2; 16824: data <= 'd0; 16825: data <= 'd0; 16826: data <= 'd0; 16827: data <= 'd0; 16828: data <= 'd0; 16829: data <= 'd0; 16830: data <= 'd0; 16831: data <= 'd0; 16832: data <= 'd0; 16833: data <= 'd0; 16834: data <= 'd0; 16835: data <= 'd0; 16836: data <= 'd0; 16837: data <= 'd0; 16838: data <= 'd0; 16839: data <= 'd0; 16840: data <= 'd2; 16841: data <= 'd5; 16842: data <= 'd3; 16843: data <= 'd6; 16844: data <= 'd3; 16845: data <= 'd1; 16846: data <= 'd1; 16847: data <= 'd1; 16848: data <= 'd1; 16849: data <= 'd1; 16850: data <= 'd1; 16851: data <= 'd1; 16852: data <= 'd1; 16853: data <= 'd1; 16854: data <= 'd3; 16855: data <= 'd2; 16856: data <= 'd0; 16857: data <= 'd0; 16858: data <= 'd0; 16859: data <= 'd0; 16860: data <= 'd0; 16861: data <= 'd0; 16862: data <= 'd0; 16863: data <= 'd0; 16864: data <= 'd0; 16865: data <= 'd0; 16866: data <= 'd0; 16867: data <= 'd0; 16868: data <= 'd0; 16869: data <= 'd0; 16870: data <= 'd0; 16871: data <= 'd0; 16872: data <= 'd2; 16873: data <= 'd5; 16874: data <= 'd3; 16875: data <= 'd1; 16876: data <= 'd1; 16877: data <= 'd1; 16878: data <= 'd5; 16879: data <= 'd5; 16880: data <= 'd5; 16881: data <= 'd5; 16882: data <= 'd5; 16883: data <= 'd5; 16884: data <= 'd5; 16885: data <= 'd1; 16886: data <= 'd1; 16887: data <= 'd2; 16888: data <= 'd0; 16889: data <= 'd0; 16890: data <= 'd0; 16891: data <= 'd0; 16892: data <= 'd0; 16893: data <= 'd0; 16894: data <= 'd0; 16895: data <= 'd0; 16896: data <= 'd0; 16897: data <= 'd0; 16898: data <= 'd0; 16899: data <= 'd0; 16900: data <= 'd0; 16901: data <= 'd0; 16902: data <= 'd0; 16903: data <= 'd0; 16904: data <= 'd2; 16905: data <= 'd6; 16906: data <= 'd1; 16907: data <= 'd5; 16908: data <= 'd2; 16909: data <= 'd2; 16910: data <= 'd2; 16911: data <= 'd2; 16912: data <= 'd2; 16913: data <= 'd2; 16914: data <= 'd2; 16915: data <= 'd2; 16916: data <= 'd2; 16917: data <= 'd2; 16918: data <= 'd5; 16919: data <= 'd2; 16920: data <= 'd0; 16921: data <= 'd0; 16922: data <= 'd0; 16923: data <= 'd0; 16924: data <= 'd0; 16925: data <= 'd0; 16926: data <= 'd0; 16927: data <= 'd0; 16928: data <= 'd0; 16929: data <= 'd0; 16930: data <= 'd0; 16931: data <= 'd0; 16932: data <= 'd0; 16933: data <= 'd0; 16934: data <= 'd2; 16935: data <= 'd2; 16936: data <= 'd5; 16937: data <= 'd6; 16938: data <= 'd5; 16939: data <= 'd2; 16940: data <= 'd8; 16941: data <= 'd8; 16942: data <= 'd8; 16943: data <= 'd8; 16944: data <= 'd8; 16945: data <= 'd9; 16946: data <= 'd9; 16947: data <= 'd8; 16948: data <= 'd8; 16949: data <= 'd8; 16950: data <= 'd2; 16951: data <= 'd2; 16952: data <= 'd0; 16953: data <= 'd0; 16954: data <= 'd0; 16955: data <= 'd0; 16956: data <= 'd0; 16957: data <= 'd0; 16958: data <= 'd0; 16959: data <= 'd0; 16960: data <= 'd0; 16961: data <= 'd0; 16962: data <= 'd0; 16963: data <= 'd0; 16964: data <= 'd0; 16965: data <= 'd0; 16966: data <= 'd2; 16967: data <= 'd3; 16968: data <= 'd6; 16969: data <= 'd3; 16970: data <= 'd2; 16971: data <= 'd8; 16972: data <= 'd8; 16973: data <= 'd9; 16974: data <= 'd9; 16975: data <= 'd10; 16976: data <= 'd2; 16977: data <= 'd9; 16978: data <= 'd11; 16979: data <= 'd10; 16980: data <= 'd2; 16981: data <= 'd9; 16982: data <= 'd2; 16983: data <= 'd2; 16984: data <= 'd0; 16985: data <= 'd0; 16986: data <= 'd0; 16987: data <= 'd0; 16988: data <= 'd0; 16989: data <= 'd0; 16990: data <= 'd0; 16991: data <= 'd0; 16992: data <= 'd0; 16993: data <= 'd0; 16994: data <= 'd0; 16995: data <= 'd0; 16996: data <= 'd0; 16997: data <= 'd0; 16998: data <= 'd2; 16999: data <= 'd1; 17000: data <= 'd3; 17001: data <= 'd1; 17002: data <= 'd2; 17003: data <= 'd10; 17004: data <= 'd10; 17005: data <= 'd9; 17006: data <= 'd10; 17007: data <= 'd10; 17008: data <= 'd11; 17009: data <= 'd10; 17010: data <= 'd11; 17011: data <= 'd11; 17012: data <= 'd10; 17013: data <= 'd10; 17014: data <= 'd2; 17015: data <= 'd0; 17016: data <= 'd0; 17017: data <= 'd0; 17018: data <= 'd0; 17019: data <= 'd0; 17020: data <= 'd0; 17021: data <= 'd0; 17022: data <= 'd0; 17023: data <= 'd0; 17024: data <= 'd0; 17025: data <= 'd0; 17026: data <= 'd0; 17027: data <= 'd0; 17028: data <= 'd0; 17029: data <= 'd0; 17030: data <= 'd0; 17031: data <= 'd2; 17032: data <= 'd1; 17033: data <= 'd5; 17034: data <= 'd2; 17035: data <= 'd8; 17036: data <= 'd9; 17037: data <= 'd9; 17038: data <= 'd10; 17039: data <= 'd10; 17040: data <= 'd10; 17041: data <= 'd10; 17042: data <= 'd8; 17043: data <= 'd8; 17044: data <= 'd10; 17045: data <= 'd9; 17046: data <= 'd2; 17047: data <= 'd0; 17048: data <= 'd0; 17049: data <= 'd0; 17050: data <= 'd0; 17051: data <= 'd0; 17052: data <= 'd0; 17053: data <= 'd0; 17054: data <= 'd0; 17055: data <= 'd0; 17056: data <= 'd0; 17057: data <= 'd0; 17058: data <= 'd0; 17059: data <= 'd0; 17060: data <= 'd0; 17061: data <= 'd0; 17062: data <= 'd0; 17063: data <= 'd0; 17064: data <= 'd2; 17065: data <= 'd2; 17066: data <= 'd2; 17067: data <= 'd8; 17068: data <= 'd8; 17069: data <= 'd9; 17070: data <= 'd9; 17071: data <= 'd10; 17072: data <= 'd10; 17073: data <= 'd10; 17074: data <= 'd9; 17075: data <= 'd9; 17076: data <= 'd10; 17077: data <= 'd9; 17078: data <= 'd2; 17079: data <= 'd0; 17080: data <= 'd0; 17081: data <= 'd0; 17082: data <= 'd0; 17083: data <= 'd0; 17084: data <= 'd0; 17085: data <= 'd0; 17086: data <= 'd0; 17087: data <= 'd0; 17088: data <= 'd0; 17089: data <= 'd0; 17090: data <= 'd0; 17091: data <= 'd0; 17092: data <= 'd0; 17093: data <= 'd0; 17094: data <= 'd0; 17095: data <= 'd0; 17096: data <= 'd0; 17097: data <= 'd0; 17098: data <= 'd0; 17099: data <= 'd2; 17100: data <= 'd5; 17101: data <= 'd5; 17102: data <= 'd8; 17103: data <= 'd9; 17104: data <= 'd9; 17105: data <= 'd9; 17106: data <= 'd9; 17107: data <= 'd9; 17108: data <= 'd9; 17109: data <= 'd2; 17110: data <= 'd0; 17111: data <= 'd0; 17112: data <= 'd0; 17113: data <= 'd0; 17114: data <= 'd0; 17115: data <= 'd0; 17116: data <= 'd0; 17117: data <= 'd0; 17118: data <= 'd0; 17119: data <= 'd0; 17120: data <= 'd0; 17121: data <= 'd0; 17122: data <= 'd0; 17123: data <= 'd0; 17124: data <= 'd0; 17125: data <= 'd0; 17126: data <= 'd0; 17127: data <= 'd0; 17128: data <= 'd0; 17129: data <= 'd0; 17130: data <= 'd2; 17131: data <= 'd7; 17132: data <= 'd1; 17133: data <= 'd1; 17134: data <= 'd1; 17135: data <= 'd3; 17136: data <= 'd3; 17137: data <= 'd3; 17138: data <= 'd5; 17139: data <= 'd5; 17140: data <= 'd3; 17141: data <= 'd1; 17142: data <= 'd2; 17143: data <= 'd0; 17144: data <= 'd0; 17145: data <= 'd0; 17146: data <= 'd0; 17147: data <= 'd0; 17148: data <= 'd0; 17149: data <= 'd0; 17150: data <= 'd0; 17151: data <= 'd0; 17152: data <= 'd0; 17153: data <= 'd0; 17154: data <= 'd0; 17155: data <= 'd0; 17156: data <= 'd0; 17157: data <= 'd0; 17158: data <= 'd0; 17159: data <= 'd0; 17160: data <= 'd0; 17161: data <= 'd2; 17162: data <= 'd7; 17163: data <= 'd7; 17164: data <= 'd7; 17165: data <= 'd1; 17166: data <= 'd1; 17167: data <= 'd3; 17168: data <= 'd3; 17169: data <= 'd3; 17170: data <= 'd1; 17171: data <= 'd1; 17172: data <= 'd3; 17173: data <= 'd1; 17174: data <= 'd2; 17175: data <= 'd2; 17176: data <= 'd0; 17177: data <= 'd0; 17178: data <= 'd0; 17179: data <= 'd0; 17180: data <= 'd0; 17181: data <= 'd0; 17182: data <= 'd0; 17183: data <= 'd0; 17184: data <= 'd0; 17185: data <= 'd0; 17186: data <= 'd0; 17187: data <= 'd0; 17188: data <= 'd0; 17189: data <= 'd0; 17190: data <= 'd0; 17191: data <= 'd0; 17192: data <= 'd2; 17193: data <= 'd8; 17194: data <= 'd10; 17195: data <= 'd10; 17196: data <= 'd5; 17197: data <= 'd1; 17198: data <= 'd1; 17199: data <= 'd1; 17200: data <= 'd3; 17201: data <= 'd3; 17202: data <= 'd1; 17203: data <= 'd1; 17204: data <= 'd1; 17205: data <= 'd1; 17206: data <= 'd8; 17207: data <= 'd9; 17208: data <= 'd2; 17209: data <= 'd0; 17210: data <= 'd0; 17211: data <= 'd0; 17212: data <= 'd0; 17213: data <= 'd0; 17214: data <= 'd0; 17215: data <= 'd0; 17216: data <= 'd0; 17217: data <= 'd0; 17218: data <= 'd0; 17219: data <= 'd0; 17220: data <= 'd0; 17221: data <= 'd0; 17222: data <= 'd0; 17223: data <= 'd0; 17224: data <= 'd2; 17225: data <= 'd9; 17226: data <= 'd10; 17227: data <= 'd9; 17228: data <= 'd2; 17229: data <= 'd2; 17230: data <= 'd2; 17231: data <= 'd2; 17232: data <= 'd2; 17233: data <= 'd5; 17234: data <= 'd5; 17235: data <= 'd5; 17236: data <= 'd2; 17237: data <= 'd2; 17238: data <= 'd8; 17239: data <= 'd9; 17240: data <= 'd2; 17241: data <= 'd0; 17242: data <= 'd0; 17243: data <= 'd0; 17244: data <= 'd0; 17245: data <= 'd0; 17246: data <= 'd0; 17247: data <= 'd0; 17248: data <= 'd0; 17249: data <= 'd0; 17250: data <= 'd0; 17251: data <= 'd0; 17252: data <= 'd0; 17253: data <= 'd0; 17254: data <= 'd0; 17255: data <= 'd0; 17256: data <= 'd0; 17257: data <= 'd2; 17258: data <= 'd2; 17259: data <= 'd2; 17260: data <= 'd2; 17261: data <= 'd1; 17262: data <= 'd1; 17263: data <= 'd3; 17264: data <= 'd3; 17265: data <= 'd3; 17266: data <= 'd1; 17267: data <= 'd3; 17268: data <= 'd3; 17269: data <= 'd2; 17270: data <= 'd2; 17271: data <= 'd2; 17272: data <= 'd0; 17273: data <= 'd0; 17274: data <= 'd0; 17275: data <= 'd0; 17276: data <= 'd0; 17277: data <= 'd0; 17278: data <= 'd0; 17279: data <= 'd0; 17280: data <= 'd0; 17281: data <= 'd0; 17282: data <= 'd0; 17283: data <= 'd0; 17284: data <= 'd0; 17285: data <= 'd0; 17286: data <= 'd0; 17287: data <= 'd0; 17288: data <= 'd0; 17289: data <= 'd0; 17290: data <= 'd0; 17291: data <= 'd0; 17292: data <= 'd2; 17293: data <= 'd4; 17294: data <= 'd7; 17295: data <= 'd7; 17296: data <= 'd4; 17297: data <= 'd2; 17298: data <= 'd5; 17299: data <= 'd4; 17300: data <= 'd2; 17301: data <= 'd0; 17302: data <= 'd0; 17303: data <= 'd0; 17304: data <= 'd0; 17305: data <= 'd0; 17306: data <= 'd0; 17307: data <= 'd0; 17308: data <= 'd0; 17309: data <= 'd0; 17310: data <= 'd0; 17311: data <= 'd0; 17312: data <= 'd0; 17313: data <= 'd0; 17314: data <= 'd0; 17315: data <= 'd0; 17316: data <= 'd0; 17317: data <= 'd0; 17318: data <= 'd0; 17319: data <= 'd0; 17320: data <= 'd0; 17321: data <= 'd0; 17322: data <= 'd0; 17323: data <= 'd0; 17324: data <= 'd0; 17325: data <= 'd2; 17326: data <= 'd4; 17327: data <= 'd7; 17328: data <= 'd2; 17329: data <= 'd4; 17330: data <= 'd4; 17331: data <= 'd2; 17332: data <= 'd0; 17333: data <= 'd0; 17334: data <= 'd0; 17335: data <= 'd0; 17336: data <= 'd0; 17337: data <= 'd0; 17338: data <= 'd0; 17339: data <= 'd0; 17340: data <= 'd0; 17341: data <= 'd0; 17342: data <= 'd0; 17343: data <= 'd0; 17344: data <= 'd0; 17345: data <= 'd0; 17346: data <= 'd0; 17347: data <= 'd0; 17348: data <= 'd0; 17349: data <= 'd0; 17350: data <= 'd0; 17351: data <= 'd0; 17352: data <= 'd0; 17353: data <= 'd0; 17354: data <= 'd0; 17355: data <= 'd0; 17356: data <= 'd0; 17357: data <= 'd0; 17358: data <= 'd2; 17359: data <= 'd2; 17360: data <= 'd2; 17361: data <= 'd2; 17362: data <= 'd2; 17363: data <= 'd0; 17364: data <= 'd0; 17365: data <= 'd0; 17366: data <= 'd0; 17367: data <= 'd0; 17368: data <= 'd0; 17369: data <= 'd0; 17370: data <= 'd0; 17371: data <= 'd0; 17372: data <= 'd0; 17373: data <= 'd0; 17374: data <= 'd0; 17375: data <= 'd0; 17376: data <= 'd0; 17377: data <= 'd0; 17378: data <= 'd0; 17379: data <= 'd0; 17380: data <= 'd0; 17381: data <= 'd0; 17382: data <= 'd0; 17383: data <= 'd0; 17384: data <= 'd0; 17385: data <= 'd0; 17386: data <= 'd0; 17387: data <= 'd0; 17388: data <= 'd0; 17389: data <= 'd0; 17390: data <= 'd0; 17391: data <= 'd0; 17392: data <= 'd0; 17393: data <= 'd0; 17394: data <= 'd0; 17395: data <= 'd0; 17396: data <= 'd0; 17397: data <= 'd0; 17398: data <= 'd0; 17399: data <= 'd0; 17400: data <= 'd0; 17401: data <= 'd0; 17402: data <= 'd0; 17403: data <= 'd0; 17404: data <= 'd0; 17405: data <= 'd0; 17406: data <= 'd0; 17407: data <= 'd0; 17408: data <= 'd0; 17409: data <= 'd0; 17410: data <= 'd0; 17411: data <= 'd0; 17412: data <= 'd0; 17413: data <= 'd0; 17414: data <= 'd0; 17415: data <= 'd0; 17416: data <= 'd0; 17417: data <= 'd0; 17418: data <= 'd0; 17419: data <= 'd0; 17420: data <= 'd0; 17421: data <= 'd0; 17422: data <= 'd0; 17423: data <= 'd0; 17424: data <= 'd0; 17425: data <= 'd0; 17426: data <= 'd0; 17427: data <= 'd0; 17428: data <= 'd0; 17429: data <= 'd0; 17430: data <= 'd0; 17431: data <= 'd0; 17432: data <= 'd0; 17433: data <= 'd0; 17434: data <= 'd0; 17435: data <= 'd0; 17436: data <= 'd0; 17437: data <= 'd0; 17438: data <= 'd0; 17439: data <= 'd0; 17440: data <= 'd0; 17441: data <= 'd0; 17442: data <= 'd0; 17443: data <= 'd0; 17444: data <= 'd0; 17445: data <= 'd0; 17446: data <= 'd0; 17447: data <= 'd0; 17448: data <= 'd0; 17449: data <= 'd0; 17450: data <= 'd0; 17451: data <= 'd0; 17452: data <= 'd0; 17453: data <= 'd0; 17454: data <= 'd0; 17455: data <= 'd0; 17456: data <= 'd0; 17457: data <= 'd0; 17458: data <= 'd0; 17459: data <= 'd0; 17460: data <= 'd0; 17461: data <= 'd0; 17462: data <= 'd0; 17463: data <= 'd0; 17464: data <= 'd0; 17465: data <= 'd0; 17466: data <= 'd0; 17467: data <= 'd0; 17468: data <= 'd0; 17469: data <= 'd0; 17470: data <= 'd0; 17471: data <= 'd0; 17472: data <= 'd0; 17473: data <= 'd0; 17474: data <= 'd0; 17475: data <= 'd0; 17476: data <= 'd0; 17477: data <= 'd0; 17478: data <= 'd0; 17479: data <= 'd0; 17480: data <= 'd0; 17481: data <= 'd0; 17482: data <= 'd0; 17483: data <= 'd0; 17484: data <= 'd0; 17485: data <= 'd0; 17486: data <= 'd0; 17487: data <= 'd0; 17488: data <= 'd0; 17489: data <= 'd0; 17490: data <= 'd0; 17491: data <= 'd0; 17492: data <= 'd0; 17493: data <= 'd0; 17494: data <= 'd0; 17495: data <= 'd0; 17496: data <= 'd0; 17497: data <= 'd0; 17498: data <= 'd0; 17499: data <= 'd0; 17500: data <= 'd0; 17501: data <= 'd0; 17502: data <= 'd0; 17503: data <= 'd0; 17504: data <= 'd0; 17505: data <= 'd0; 17506: data <= 'd0; 17507: data <= 'd0; 17508: data <= 'd0; 17509: data <= 'd0; 17510: data <= 'd0; 17511: data <= 'd0; 17512: data <= 'd0; 17513: data <= 'd0; 17514: data <= 'd0; 17515: data <= 'd0; 17516: data <= 'd0; 17517: data <= 'd0; 17518: data <= 'd0; 17519: data <= 'd0; 17520: data <= 'd0; 17521: data <= 'd0; 17522: data <= 'd0; 17523: data <= 'd0; 17524: data <= 'd0; 17525: data <= 'd0; 17526: data <= 'd0; 17527: data <= 'd0; 17528: data <= 'd0; 17529: data <= 'd0; 17530: data <= 'd0; 17531: data <= 'd0; 17532: data <= 'd0; 17533: data <= 'd0; 17534: data <= 'd0; 17535: data <= 'd0; 17536: data <= 'd0; 17537: data <= 'd0; 17538: data <= 'd0; 17539: data <= 'd0; 17540: data <= 'd0; 17541: data <= 'd0; 17542: data <= 'd0; 17543: data <= 'd0; 17544: data <= 'd0; 17545: data <= 'd0; 17546: data <= 'd0; 17547: data <= 'd0; 17548: data <= 'd0; 17549: data <= 'd0; 17550: data <= 'd0; 17551: data <= 'd0; 17552: data <= 'd0; 17553: data <= 'd0; 17554: data <= 'd0; 17555: data <= 'd0; 17556: data <= 'd0; 17557: data <= 'd0; 17558: data <= 'd0; 17559: data <= 'd0; 17560: data <= 'd0; 17561: data <= 'd0; 17562: data <= 'd0; 17563: data <= 'd0; 17564: data <= 'd0; 17565: data <= 'd0; 17566: data <= 'd0; 17567: data <= 'd0; 17568: data <= 'd0; 17569: data <= 'd0; 17570: data <= 'd0; 17571: data <= 'd0; 17572: data <= 'd0; 17573: data <= 'd0; 17574: data <= 'd0; 17575: data <= 'd0; 17576: data <= 'd0; 17577: data <= 'd0; 17578: data <= 'd0; 17579: data <= 'd0; 17580: data <= 'd0; 17581: data <= 'd0; 17582: data <= 'd0; 17583: data <= 'd0; 17584: data <= 'd0; 17585: data <= 'd0; 17586: data <= 'd0; 17587: data <= 'd0; 17588: data <= 'd0; 17589: data <= 'd0; 17590: data <= 'd0; 17591: data <= 'd0; 17592: data <= 'd0; 17593: data <= 'd0; 17594: data <= 'd0; 17595: data <= 'd0; 17596: data <= 'd0; 17597: data <= 'd0; 17598: data <= 'd0; 17599: data <= 'd0; 17600: data <= 'd0; 17601: data <= 'd0; 17602: data <= 'd0; 17603: data <= 'd0; 17604: data <= 'd0; 17605: data <= 'd0; 17606: data <= 'd0; 17607: data <= 'd0; 17608: data <= 'd0; 17609: data <= 'd0; 17610: data <= 'd0; 17611: data <= 'd0; 17612: data <= 'd0; 17613: data <= 'd0; 17614: data <= 'd0; 17615: data <= 'd0; 17616: data <= 'd0; 17617: data <= 'd0; 17618: data <= 'd0; 17619: data <= 'd0; 17620: data <= 'd0; 17621: data <= 'd0; 17622: data <= 'd0; 17623: data <= 'd0; 17624: data <= 'd0; 17625: data <= 'd0; 17626: data <= 'd0; 17627: data <= 'd0; 17628: data <= 'd0; 17629: data <= 'd0; 17630: data <= 'd0; 17631: data <= 'd0; 17632: data <= 'd0; 17633: data <= 'd0; 17634: data <= 'd0; 17635: data <= 'd0; 17636: data <= 'd0; 17637: data <= 'd0; 17638: data <= 'd0; 17639: data <= 'd0; 17640: data <= 'd0; 17641: data <= 'd0; 17642: data <= 'd0; 17643: data <= 'd0; 17644: data <= 'd0; 17645: data <= 'd0; 17646: data <= 'd0; 17647: data <= 'd0; 17648: data <= 'd0; 17649: data <= 'd0; 17650: data <= 'd0; 17651: data <= 'd0; 17652: data <= 'd0; 17653: data <= 'd0; 17654: data <= 'd0; 17655: data <= 'd0; 17656: data <= 'd0; 17657: data <= 'd0; 17658: data <= 'd0; 17659: data <= 'd0; 17660: data <= 'd0; 17661: data <= 'd0; 17662: data <= 'd0; 17663: data <= 'd0; 17664: data <= 'd0; 17665: data <= 'd0; 17666: data <= 'd0; 17667: data <= 'd0; 17668: data <= 'd0; 17669: data <= 'd0; 17670: data <= 'd0; 17671: data <= 'd0; 17672: data <= 'd0; 17673: data <= 'd0; 17674: data <= 'd0; 17675: data <= 'd0; 17676: data <= 'd0; 17677: data <= 'd0; 17678: data <= 'd0; 17679: data <= 'd0; 17680: data <= 'd0; 17681: data <= 'd0; 17682: data <= 'd0; 17683: data <= 'd0; 17684: data <= 'd0; 17685: data <= 'd0; 17686: data <= 'd0; 17687: data <= 'd0; 17688: data <= 'd0; 17689: data <= 'd0; 17690: data <= 'd0; 17691: data <= 'd0; 17692: data <= 'd0; 17693: data <= 'd0; 17694: data <= 'd0; 17695: data <= 'd0; 17696: data <= 'd0; 17697: data <= 'd0; 17698: data <= 'd0; 17699: data <= 'd0; 17700: data <= 'd0; 17701: data <= 'd0; 17702: data <= 'd0; 17703: data <= 'd0; 17704: data <= 'd0; 17705: data <= 'd0; 17706: data <= 'd0; 17707: data <= 'd0; 17708: data <= 'd0; 17709: data <= 'd2; 17710: data <= 'd2; 17711: data <= 'd2; 17712: data <= 'd2; 17713: data <= 'd2; 17714: data <= 'd2; 17715: data <= 'd0; 17716: data <= 'd0; 17717: data <= 'd0; 17718: data <= 'd0; 17719: data <= 'd0; 17720: data <= 'd0; 17721: data <= 'd0; 17722: data <= 'd0; 17723: data <= 'd0; 17724: data <= 'd0; 17725: data <= 'd0; 17726: data <= 'd0; 17727: data <= 'd0; 17728: data <= 'd0; 17729: data <= 'd0; 17730: data <= 'd0; 17731: data <= 'd0; 17732: data <= 'd0; 17733: data <= 'd0; 17734: data <= 'd0; 17735: data <= 'd0; 17736: data <= 'd0; 17737: data <= 'd0; 17738: data <= 'd0; 17739: data <= 'd2; 17740: data <= 'd2; 17741: data <= 'd6; 17742: data <= 'd6; 17743: data <= 'd6; 17744: data <= 'd6; 17745: data <= 'd6; 17746: data <= 'd6; 17747: data <= 'd2; 17748: data <= 'd2; 17749: data <= 'd0; 17750: data <= 'd0; 17751: data <= 'd0; 17752: data <= 'd0; 17753: data <= 'd0; 17754: data <= 'd0; 17755: data <= 'd0; 17756: data <= 'd0; 17757: data <= 'd0; 17758: data <= 'd0; 17759: data <= 'd0; 17760: data <= 'd0; 17761: data <= 'd0; 17762: data <= 'd0; 17763: data <= 'd0; 17764: data <= 'd0; 17765: data <= 'd0; 17766: data <= 'd0; 17767: data <= 'd0; 17768: data <= 'd0; 17769: data <= 'd0; 17770: data <= 'd2; 17771: data <= 'd1; 17772: data <= 'd3; 17773: data <= 'd6; 17774: data <= 'd6; 17775: data <= 'd6; 17776: data <= 'd6; 17777: data <= 'd6; 17778: data <= 'd6; 17779: data <= 'd6; 17780: data <= 'd3; 17781: data <= 'd2; 17782: data <= 'd0; 17783: data <= 'd0; 17784: data <= 'd0; 17785: data <= 'd0; 17786: data <= 'd0; 17787: data <= 'd0; 17788: data <= 'd0; 17789: data <= 'd0; 17790: data <= 'd0; 17791: data <= 'd0; 17792: data <= 'd0; 17793: data <= 'd0; 17794: data <= 'd0; 17795: data <= 'd0; 17796: data <= 'd0; 17797: data <= 'd0; 17798: data <= 'd0; 17799: data <= 'd0; 17800: data <= 'd0; 17801: data <= 'd2; 17802: data <= 'd1; 17803: data <= 'd1; 17804: data <= 'd1; 17805: data <= 'd3; 17806: data <= 'd6; 17807: data <= 'd6; 17808: data <= 'd6; 17809: data <= 'd6; 17810: data <= 'd6; 17811: data <= 'd3; 17812: data <= 'd1; 17813: data <= 'd1; 17814: data <= 'd2; 17815: data <= 'd0; 17816: data <= 'd0; 17817: data <= 'd0; 17818: data <= 'd0; 17819: data <= 'd0; 17820: data <= 'd0; 17821: data <= 'd0; 17822: data <= 'd0; 17823: data <= 'd0; 17824: data <= 'd0; 17825: data <= 'd0; 17826: data <= 'd0; 17827: data <= 'd0; 17828: data <= 'd0; 17829: data <= 'd0; 17830: data <= 'd0; 17831: data <= 'd0; 17832: data <= 'd0; 17833: data <= 'd2; 17834: data <= 'd1; 17835: data <= 'd1; 17836: data <= 'd5; 17837: data <= 'd5; 17838: data <= 'd5; 17839: data <= 'd1; 17840: data <= 'd1; 17841: data <= 'd1; 17842: data <= 'd1; 17843: data <= 'd1; 17844: data <= 'd5; 17845: data <= 'd5; 17846: data <= 'd2; 17847: data <= 'd0; 17848: data <= 'd0; 17849: data <= 'd0; 17850: data <= 'd0; 17851: data <= 'd0; 17852: data <= 'd0; 17853: data <= 'd0; 17854: data <= 'd0; 17855: data <= 'd0; 17856: data <= 'd0; 17857: data <= 'd0; 17858: data <= 'd0; 17859: data <= 'd0; 17860: data <= 'd0; 17861: data <= 'd0; 17862: data <= 'd0; 17863: data <= 'd0; 17864: data <= 'd2; 17865: data <= 'd1; 17866: data <= 'd5; 17867: data <= 'd5; 17868: data <= 'd3; 17869: data <= 'd6; 17870: data <= 'd6; 17871: data <= 'd6; 17872: data <= 'd6; 17873: data <= 'd6; 17874: data <= 'd6; 17875: data <= 'd6; 17876: data <= 'd6; 17877: data <= 'd3; 17878: data <= 'd5; 17879: data <= 'd2; 17880: data <= 'd0; 17881: data <= 'd0; 17882: data <= 'd0; 17883: data <= 'd0; 17884: data <= 'd0; 17885: data <= 'd0; 17886: data <= 'd0; 17887: data <= 'd0; 17888: data <= 'd0; 17889: data <= 'd0; 17890: data <= 'd0; 17891: data <= 'd0; 17892: data <= 'd0; 17893: data <= 'd0; 17894: data <= 'd0; 17895: data <= 'd0; 17896: data <= 'd2; 17897: data <= 'd5; 17898: data <= 'd3; 17899: data <= 'd6; 17900: data <= 'd3; 17901: data <= 'd1; 17902: data <= 'd1; 17903: data <= 'd1; 17904: data <= 'd1; 17905: data <= 'd1; 17906: data <= 'd1; 17907: data <= 'd1; 17908: data <= 'd1; 17909: data <= 'd1; 17910: data <= 'd3; 17911: data <= 'd2; 17912: data <= 'd0; 17913: data <= 'd0; 17914: data <= 'd0; 17915: data <= 'd0; 17916: data <= 'd0; 17917: data <= 'd0; 17918: data <= 'd0; 17919: data <= 'd0; 17920: data <= 'd0; 17921: data <= 'd0; 17922: data <= 'd0; 17923: data <= 'd0; 17924: data <= 'd0; 17925: data <= 'd0; 17926: data <= 'd0; 17927: data <= 'd0; 17928: data <= 'd2; 17929: data <= 'd5; 17930: data <= 'd3; 17931: data <= 'd1; 17932: data <= 'd1; 17933: data <= 'd1; 17934: data <= 'd5; 17935: data <= 'd5; 17936: data <= 'd5; 17937: data <= 'd5; 17938: data <= 'd5; 17939: data <= 'd5; 17940: data <= 'd5; 17941: data <= 'd1; 17942: data <= 'd1; 17943: data <= 'd2; 17944: data <= 'd0; 17945: data <= 'd0; 17946: data <= 'd0; 17947: data <= 'd0; 17948: data <= 'd0; 17949: data <= 'd0; 17950: data <= 'd0; 17951: data <= 'd0; 17952: data <= 'd0; 17953: data <= 'd0; 17954: data <= 'd0; 17955: data <= 'd0; 17956: data <= 'd0; 17957: data <= 'd0; 17958: data <= 'd0; 17959: data <= 'd0; 17960: data <= 'd2; 17961: data <= 'd6; 17962: data <= 'd1; 17963: data <= 'd5; 17964: data <= 'd2; 17965: data <= 'd2; 17966: data <= 'd2; 17967: data <= 'd2; 17968: data <= 'd2; 17969: data <= 'd2; 17970: data <= 'd2; 17971: data <= 'd2; 17972: data <= 'd2; 17973: data <= 'd2; 17974: data <= 'd5; 17975: data <= 'd2; 17976: data <= 'd0; 17977: data <= 'd0; 17978: data <= 'd0; 17979: data <= 'd0; 17980: data <= 'd0; 17981: data <= 'd0; 17982: data <= 'd0; 17983: data <= 'd0; 17984: data <= 'd0; 17985: data <= 'd0; 17986: data <= 'd0; 17987: data <= 'd0; 17988: data <= 'd0; 17989: data <= 'd0; 17990: data <= 'd2; 17991: data <= 'd2; 17992: data <= 'd2; 17993: data <= 'd1; 17994: data <= 'd5; 17995: data <= 'd2; 17996: data <= 'd8; 17997: data <= 'd8; 17998: data <= 'd8; 17999: data <= 'd8; 18000: data <= 'd8; 18001: data <= 'd9; 18002: data <= 'd9; 18003: data <= 'd8; 18004: data <= 'd8; 18005: data <= 'd8; 18006: data <= 'd2; 18007: data <= 'd2; 18008: data <= 'd0; 18009: data <= 'd0; 18010: data <= 'd0; 18011: data <= 'd0; 18012: data <= 'd0; 18013: data <= 'd0; 18014: data <= 'd0; 18015: data <= 'd0; 18016: data <= 'd0; 18017: data <= 'd0; 18018: data <= 'd0; 18019: data <= 'd0; 18020: data <= 'd0; 18021: data <= 'd0; 18022: data <= 'd2; 18023: data <= 'd1; 18024: data <= 'd2; 18025: data <= 'd1; 18026: data <= 'd2; 18027: data <= 'd8; 18028: data <= 'd8; 18029: data <= 'd9; 18030: data <= 'd9; 18031: data <= 'd2; 18032: data <= 'd9; 18033: data <= 'd11; 18034: data <= 'd11; 18035: data <= 'd10; 18036: data <= 'd2; 18037: data <= 'd9; 18038: data <= 'd2; 18039: data <= 'd2; 18040: data <= 'd0; 18041: data <= 'd0; 18042: data <= 'd0; 18043: data <= 'd0; 18044: data <= 'd0; 18045: data <= 'd0; 18046: data <= 'd0; 18047: data <= 'd0; 18048: data <= 'd0; 18049: data <= 'd0; 18050: data <= 'd0; 18051: data <= 'd0; 18052: data <= 'd0; 18053: data <= 'd0; 18054: data <= 'd2; 18055: data <= 'd5; 18056: data <= 'd1; 18057: data <= 'd2; 18058: data <= 'd9; 18059: data <= 'd10; 18060: data <= 'd9; 18061: data <= 'd9; 18062: data <= 'd10; 18063: data <= 'd11; 18064: data <= 'd10; 18065: data <= 'd11; 18066: data <= 'd11; 18067: data <= 'd10; 18068: data <= 'd11; 18069: data <= 'd10; 18070: data <= 'd9; 18071: data <= 'd2; 18072: data <= 'd0; 18073: data <= 'd0; 18074: data <= 'd0; 18075: data <= 'd0; 18076: data <= 'd0; 18077: data <= 'd0; 18078: data <= 'd0; 18079: data <= 'd0; 18080: data <= 'd0; 18081: data <= 'd0; 18082: data <= 'd0; 18083: data <= 'd0; 18084: data <= 'd0; 18085: data <= 'd0; 18086: data <= 'd0; 18087: data <= 'd2; 18088: data <= 'd5; 18089: data <= 'd5; 18090: data <= 'd2; 18091: data <= 'd8; 18092: data <= 'd9; 18093: data <= 'd9; 18094: data <= 'd10; 18095: data <= 'd10; 18096: data <= 'd10; 18097: data <= 'd8; 18098: data <= 'd8; 18099: data <= 'd10; 18100: data <= 'd10; 18101: data <= 'd9; 18102: data <= 'd2; 18103: data <= 'd0; 18104: data <= 'd0; 18105: data <= 'd0; 18106: data <= 'd0; 18107: data <= 'd0; 18108: data <= 'd0; 18109: data <= 'd0; 18110: data <= 'd0; 18111: data <= 'd0; 18112: data <= 'd0; 18113: data <= 'd0; 18114: data <= 'd0; 18115: data <= 'd0; 18116: data <= 'd0; 18117: data <= 'd0; 18118: data <= 'd0; 18119: data <= 'd0; 18120: data <= 'd2; 18121: data <= 'd2; 18122: data <= 'd2; 18123: data <= 'd8; 18124: data <= 'd8; 18125: data <= 'd9; 18126: data <= 'd9; 18127: data <= 'd10; 18128: data <= 'd10; 18129: data <= 'd9; 18130: data <= 'd9; 18131: data <= 'd10; 18132: data <= 'd10; 18133: data <= 'd9; 18134: data <= 'd2; 18135: data <= 'd0; 18136: data <= 'd0; 18137: data <= 'd0; 18138: data <= 'd0; 18139: data <= 'd0; 18140: data <= 'd0; 18141: data <= 'd0; 18142: data <= 'd0; 18143: data <= 'd0; 18144: data <= 'd0; 18145: data <= 'd0; 18146: data <= 'd0; 18147: data <= 'd0; 18148: data <= 'd0; 18149: data <= 'd0; 18150: data <= 'd0; 18151: data <= 'd0; 18152: data <= 'd0; 18153: data <= 'd0; 18154: data <= 'd2; 18155: data <= 'd2; 18156: data <= 'd5; 18157: data <= 'd5; 18158: data <= 'd8; 18159: data <= 'd9; 18160: data <= 'd9; 18161: data <= 'd9; 18162: data <= 'd9; 18163: data <= 'd9; 18164: data <= 'd9; 18165: data <= 'd5; 18166: data <= 'd2; 18167: data <= 'd0; 18168: data <= 'd0; 18169: data <= 'd0; 18170: data <= 'd0; 18171: data <= 'd0; 18172: data <= 'd0; 18173: data <= 'd0; 18174: data <= 'd0; 18175: data <= 'd0; 18176: data <= 'd0; 18177: data <= 'd0; 18178: data <= 'd0; 18179: data <= 'd0; 18180: data <= 'd0; 18181: data <= 'd0; 18182: data <= 'd0; 18183: data <= 'd0; 18184: data <= 'd0; 18185: data <= 'd2; 18186: data <= 'd7; 18187: data <= 'd1; 18188: data <= 'd1; 18189: data <= 'd1; 18190: data <= 'd3; 18191: data <= 'd3; 18192: data <= 'd3; 18193: data <= 'd5; 18194: data <= 'd5; 18195: data <= 'd3; 18196: data <= 'd3; 18197: data <= 'd1; 18198: data <= 'd2; 18199: data <= 'd0; 18200: data <= 'd0; 18201: data <= 'd0; 18202: data <= 'd0; 18203: data <= 'd0; 18204: data <= 'd0; 18205: data <= 'd0; 18206: data <= 'd0; 18207: data <= 'd0; 18208: data <= 'd0; 18209: data <= 'd0; 18210: data <= 'd0; 18211: data <= 'd0; 18212: data <= 'd0; 18213: data <= 'd0; 18214: data <= 'd0; 18215: data <= 'd0; 18216: data <= 'd0; 18217: data <= 'd2; 18218: data <= 'd7; 18219: data <= 'd7; 18220: data <= 'd1; 18221: data <= 'd1; 18222: data <= 'd3; 18223: data <= 'd3; 18224: data <= 'd3; 18225: data <= 'd1; 18226: data <= 'd1; 18227: data <= 'd3; 18228: data <= 'd3; 18229: data <= 'd1; 18230: data <= 'd2; 18231: data <= 'd0; 18232: data <= 'd0; 18233: data <= 'd0; 18234: data <= 'd0; 18235: data <= 'd0; 18236: data <= 'd0; 18237: data <= 'd0; 18238: data <= 'd0; 18239: data <= 'd0; 18240: data <= 'd0; 18241: data <= 'd0; 18242: data <= 'd0; 18243: data <= 'd0; 18244: data <= 'd0; 18245: data <= 'd0; 18246: data <= 'd0; 18247: data <= 'd0; 18248: data <= 'd2; 18249: data <= 'd9; 18250: data <= 'd9; 18251: data <= 'd7; 18252: data <= 'd1; 18253: data <= 'd1; 18254: data <= 'd1; 18255: data <= 'd3; 18256: data <= 'd3; 18257: data <= 'd1; 18258: data <= 'd1; 18259: data <= 'd3; 18260: data <= 'd1; 18261: data <= 'd1; 18262: data <= 'd8; 18263: data <= 'd2; 18264: data <= 'd0; 18265: data <= 'd0; 18266: data <= 'd0; 18267: data <= 'd0; 18268: data <= 'd0; 18269: data <= 'd0; 18270: data <= 'd0; 18271: data <= 'd0; 18272: data <= 'd0; 18273: data <= 'd0; 18274: data <= 'd0; 18275: data <= 'd0; 18276: data <= 'd0; 18277: data <= 'd0; 18278: data <= 'd0; 18279: data <= 'd0; 18280: data <= 'd2; 18281: data <= 'd9; 18282: data <= 'd9; 18283: data <= 'd2; 18284: data <= 'd2; 18285: data <= 'd2; 18286: data <= 'd2; 18287: data <= 'd2; 18288: data <= 'd5; 18289: data <= 'd5; 18290: data <= 'd5; 18291: data <= 'd2; 18292: data <= 'd2; 18293: data <= 'd2; 18294: data <= 'd8; 18295: data <= 'd2; 18296: data <= 'd0; 18297: data <= 'd0; 18298: data <= 'd0; 18299: data <= 'd0; 18300: data <= 'd0; 18301: data <= 'd0; 18302: data <= 'd0; 18303: data <= 'd0; 18304: data <= 'd0; 18305: data <= 'd0; 18306: data <= 'd0; 18307: data <= 'd0; 18308: data <= 'd0; 18309: data <= 'd0; 18310: data <= 'd0; 18311: data <= 'd0; 18312: data <= 'd0; 18313: data <= 'd2; 18314: data <= 'd2; 18315: data <= 'd2; 18316: data <= 'd1; 18317: data <= 'd1; 18318: data <= 'd3; 18319: data <= 'd3; 18320: data <= 'd3; 18321: data <= 'd1; 18322: data <= 'd3; 18323: data <= 'd3; 18324: data <= 'd3; 18325: data <= 'd2; 18326: data <= 'd2; 18327: data <= 'd0; 18328: data <= 'd0; 18329: data <= 'd0; 18330: data <= 'd0; 18331: data <= 'd0; 18332: data <= 'd0; 18333: data <= 'd0; 18334: data <= 'd0; 18335: data <= 'd0; 18336: data <= 'd0; 18337: data <= 'd0; 18338: data <= 'd0; 18339: data <= 'd0; 18340: data <= 'd0; 18341: data <= 'd0; 18342: data <= 'd0; 18343: data <= 'd0; 18344: data <= 'd0; 18345: data <= 'd0; 18346: data <= 'd0; 18347: data <= 'd2; 18348: data <= 'd4; 18349: data <= 'd7; 18350: data <= 'd7; 18351: data <= 'd2; 18352: data <= 'd2; 18353: data <= 'd2; 18354: data <= 'd2; 18355: data <= 'd4; 18356: data <= 'd4; 18357: data <= 'd2; 18358: data <= 'd0; 18359: data <= 'd0; 18360: data <= 'd0; 18361: data <= 'd0; 18362: data <= 'd0; 18363: data <= 'd0; 18364: data <= 'd0; 18365: data <= 'd0; 18366: data <= 'd0; 18367: data <= 'd0; 18368: data <= 'd0; 18369: data <= 'd0; 18370: data <= 'd0; 18371: data <= 'd0; 18372: data <= 'd0; 18373: data <= 'd0; 18374: data <= 'd0; 18375: data <= 'd0; 18376: data <= 'd0; 18377: data <= 'd0; 18378: data <= 'd0; 18379: data <= 'd2; 18380: data <= 'd4; 18381: data <= 'd7; 18382: data <= 'd2; 18383: data <= 'd0; 18384: data <= 'd0; 18385: data <= 'd0; 18386: data <= 'd2; 18387: data <= 'd2; 18388: data <= 'd2; 18389: data <= 'd2; 18390: data <= 'd0; 18391: data <= 'd0; 18392: data <= 'd0; 18393: data <= 'd0; 18394: data <= 'd0; 18395: data <= 'd0; 18396: data <= 'd0; 18397: data <= 'd0; 18398: data <= 'd0; 18399: data <= 'd0; 18400: data <= 'd0; 18401: data <= 'd0; 18402: data <= 'd0; 18403: data <= 'd0; 18404: data <= 'd0; 18405: data <= 'd0; 18406: data <= 'd0; 18407: data <= 'd0; 18408: data <= 'd0; 18409: data <= 'd0; 18410: data <= 'd0; 18411: data <= 'd2; 18412: data <= 'd2; 18413: data <= 'd2; 18414: data <= 'd0; 18415: data <= 'd0; 18416: data <= 'd0; 18417: data <= 'd0; 18418: data <= 'd0; 18419: data <= 'd0; 18420: data <= 'd0; 18421: data <= 'd0; 18422: data <= 'd0; 18423: data <= 'd0; 18424: data <= 'd0; 18425: data <= 'd0; 18426: data <= 'd0; 18427: data <= 'd0; 18428: data <= 'd0; 18429: data <= 'd0; 18430: data <= 'd0; 18431: data <= 'd0; 18432: data <= 'd0; 18433: data <= 'd0; 18434: data <= 'd0; 18435: data <= 'd0; 18436: data <= 'd0; 18437: data <= 'd0; 18438: data <= 'd0; 18439: data <= 'd0; 18440: data <= 'd0; 18441: data <= 'd0; 18442: data <= 'd0; 18443: data <= 'd0; 18444: data <= 'd0; 18445: data <= 'd0; 18446: data <= 'd0; 18447: data <= 'd0; 18448: data <= 'd0; 18449: data <= 'd0; 18450: data <= 'd0; 18451: data <= 'd0; 18452: data <= 'd0; 18453: data <= 'd0; 18454: data <= 'd0; 18455: data <= 'd0; 18456: data <= 'd0; 18457: data <= 'd0; 18458: data <= 'd0; 18459: data <= 'd0; 18460: data <= 'd0; 18461: data <= 'd0; 18462: data <= 'd0; 18463: data <= 'd0; 18464: data <= 'd0; 18465: data <= 'd0; 18466: data <= 'd0; 18467: data <= 'd0; 18468: data <= 'd0; 18469: data <= 'd0; 18470: data <= 'd0; 18471: data <= 'd0; 18472: data <= 'd0; 18473: data <= 'd0; 18474: data <= 'd0; 18475: data <= 'd0; 18476: data <= 'd0; 18477: data <= 'd0; 18478: data <= 'd0; 18479: data <= 'd0; 18480: data <= 'd0; 18481: data <= 'd0; 18482: data <= 'd0; 18483: data <= 'd0; 18484: data <= 'd0; 18485: data <= 'd0; 18486: data <= 'd0; 18487: data <= 'd0; 18488: data <= 'd0; 18489: data <= 'd0; 18490: data <= 'd0; 18491: data <= 'd0; 18492: data <= 'd0; 18493: data <= 'd0; 18494: data <= 'd0; 18495: data <= 'd0; 18496: data <= 'd0; 18497: data <= 'd0; 18498: data <= 'd0; 18499: data <= 'd0; 18500: data <= 'd0; 18501: data <= 'd0; 18502: data <= 'd0; 18503: data <= 'd0; 18504: data <= 'd0; 18505: data <= 'd0; 18506: data <= 'd0; 18507: data <= 'd0; 18508: data <= 'd0; 18509: data <= 'd0; 18510: data <= 'd0; 18511: data <= 'd0; 18512: data <= 'd0; 18513: data <= 'd0; 18514: data <= 'd0; 18515: data <= 'd0; 18516: data <= 'd0; 18517: data <= 'd0; 18518: data <= 'd0; 18519: data <= 'd0; 18520: data <= 'd0; 18521: data <= 'd0; 18522: data <= 'd0; 18523: data <= 'd0; 18524: data <= 'd0; 18525: data <= 'd0; 18526: data <= 'd0; 18527: data <= 'd0; 18528: data <= 'd0; 18529: data <= 'd0; 18530: data <= 'd0; 18531: data <= 'd0; 18532: data <= 'd0; 18533: data <= 'd0; 18534: data <= 'd0; 18535: data <= 'd0; 18536: data <= 'd0; 18537: data <= 'd0; 18538: data <= 'd0; 18539: data <= 'd0; 18540: data <= 'd0; 18541: data <= 'd0; 18542: data <= 'd0; 18543: data <= 'd0; 18544: data <= 'd0; 18545: data <= 'd0; 18546: data <= 'd0; 18547: data <= 'd0; 18548: data <= 'd0; 18549: data <= 'd0; 18550: data <= 'd0; 18551: data <= 'd0; 18552: data <= 'd0; 18553: data <= 'd0; 18554: data <= 'd0; 18555: data <= 'd0; 18556: data <= 'd0; 18557: data <= 'd0; 18558: data <= 'd0; 18559: data <= 'd0; 18560: data <= 'd0; 18561: data <= 'd0; 18562: data <= 'd0; 18563: data <= 'd0; 18564: data <= 'd0; 18565: data <= 'd0; 18566: data <= 'd0; 18567: data <= 'd0; 18568: data <= 'd0; 18569: data <= 'd0; 18570: data <= 'd0; 18571: data <= 'd0; 18572: data <= 'd0; 18573: data <= 'd0; 18574: data <= 'd0; 18575: data <= 'd0; 18576: data <= 'd0; 18577: data <= 'd0; 18578: data <= 'd0; 18579: data <= 'd0; 18580: data <= 'd0; 18581: data <= 'd0; 18582: data <= 'd0; 18583: data <= 'd0; 18584: data <= 'd0; 18585: data <= 'd0; 18586: data <= 'd0; 18587: data <= 'd0; 18588: data <= 'd0; 18589: data <= 'd0; 18590: data <= 'd0; 18591: data <= 'd0; 18592: data <= 'd0; 18593: data <= 'd0; 18594: data <= 'd0; 18595: data <= 'd0; 18596: data <= 'd0; 18597: data <= 'd0; 18598: data <= 'd0; 18599: data <= 'd0; 18600: data <= 'd0; 18601: data <= 'd0; 18602: data <= 'd0; 18603: data <= 'd0; 18604: data <= 'd0; 18605: data <= 'd0; 18606: data <= 'd0; 18607: data <= 'd0; 18608: data <= 'd0; 18609: data <= 'd0; 18610: data <= 'd0; 18611: data <= 'd0; 18612: data <= 'd0; 18613: data <= 'd0; 18614: data <= 'd0; 18615: data <= 'd0; 18616: data <= 'd0; 18617: data <= 'd0; 18618: data <= 'd0; 18619: data <= 'd0; 18620: data <= 'd0; 18621: data <= 'd0; 18622: data <= 'd0; 18623: data <= 'd0; 18624: data <= 'd0; 18625: data <= 'd0; 18626: data <= 'd0; 18627: data <= 'd0; 18628: data <= 'd0; 18629: data <= 'd0; 18630: data <= 'd0; 18631: data <= 'd0; 18632: data <= 'd0; 18633: data <= 'd0; 18634: data <= 'd0; 18635: data <= 'd0; 18636: data <= 'd0; 18637: data <= 'd0; 18638: data <= 'd0; 18639: data <= 'd0; 18640: data <= 'd0; 18641: data <= 'd0; 18642: data <= 'd0; 18643: data <= 'd0; 18644: data <= 'd0; 18645: data <= 'd0; 18646: data <= 'd0; 18647: data <= 'd0; 18648: data <= 'd0; 18649: data <= 'd0; 18650: data <= 'd0; 18651: data <= 'd0; 18652: data <= 'd0; 18653: data <= 'd0; 18654: data <= 'd0; 18655: data <= 'd0; 18656: data <= 'd0; 18657: data <= 'd0; 18658: data <= 'd0; 18659: data <= 'd0; 18660: data <= 'd0; 18661: data <= 'd0; 18662: data <= 'd0; 18663: data <= 'd0; 18664: data <= 'd0; 18665: data <= 'd0; 18666: data <= 'd0; 18667: data <= 'd0; 18668: data <= 'd0; 18669: data <= 'd0; 18670: data <= 'd0; 18671: data <= 'd0; 18672: data <= 'd0; 18673: data <= 'd0; 18674: data <= 'd0; 18675: data <= 'd0; 18676: data <= 'd0; 18677: data <= 'd0; 18678: data <= 'd0; 18679: data <= 'd0; 18680: data <= 'd0; 18681: data <= 'd0; 18682: data <= 'd0; 18683: data <= 'd0; 18684: data <= 'd0; 18685: data <= 'd0; 18686: data <= 'd0; 18687: data <= 'd0; 18688: data <= 'd0; 18689: data <= 'd0; 18690: data <= 'd0; 18691: data <= 'd0; 18692: data <= 'd0; 18693: data <= 'd0; 18694: data <= 'd0; 18695: data <= 'd0; 18696: data <= 'd0; 18697: data <= 'd0; 18698: data <= 'd0; 18699: data <= 'd0; 18700: data <= 'd0; 18701: data <= 'd2; 18702: data <= 'd2; 18703: data <= 'd2; 18704: data <= 'd2; 18705: data <= 'd2; 18706: data <= 'd0; 18707: data <= 'd0; 18708: data <= 'd0; 18709: data <= 'd0; 18710: data <= 'd0; 18711: data <= 'd0; 18712: data <= 'd0; 18713: data <= 'd0; 18714: data <= 'd0; 18715: data <= 'd0; 18716: data <= 'd0; 18717: data <= 'd0; 18718: data <= 'd0; 18719: data <= 'd0; 18720: data <= 'd0; 18721: data <= 'd0; 18722: data <= 'd0; 18723: data <= 'd0; 18724: data <= 'd0; 18725: data <= 'd0; 18726: data <= 'd0; 18727: data <= 'd0; 18728: data <= 'd0; 18729: data <= 'd0; 18730: data <= 'd0; 18731: data <= 'd2; 18732: data <= 'd2; 18733: data <= 'd6; 18734: data <= 'd6; 18735: data <= 'd6; 18736: data <= 'd6; 18737: data <= 'd6; 18738: data <= 'd2; 18739: data <= 'd2; 18740: data <= 'd0; 18741: data <= 'd0; 18742: data <= 'd0; 18743: data <= 'd0; 18744: data <= 'd0; 18745: data <= 'd0; 18746: data <= 'd0; 18747: data <= 'd0; 18748: data <= 'd0; 18749: data <= 'd0; 18750: data <= 'd0; 18751: data <= 'd0; 18752: data <= 'd0; 18753: data <= 'd0; 18754: data <= 'd0; 18755: data <= 'd0; 18756: data <= 'd0; 18757: data <= 'd0; 18758: data <= 'd0; 18759: data <= 'd0; 18760: data <= 'd0; 18761: data <= 'd0; 18762: data <= 'd2; 18763: data <= 'd3; 18764: data <= 'd6; 18765: data <= 'd6; 18766: data <= 'd6; 18767: data <= 'd6; 18768: data <= 'd6; 18769: data <= 'd6; 18770: data <= 'd6; 18771: data <= 'd3; 18772: data <= 'd2; 18773: data <= 'd0; 18774: data <= 'd0; 18775: data <= 'd0; 18776: data <= 'd0; 18777: data <= 'd0; 18778: data <= 'd0; 18779: data <= 'd0; 18780: data <= 'd0; 18781: data <= 'd0; 18782: data <= 'd0; 18783: data <= 'd0; 18784: data <= 'd0; 18785: data <= 'd0; 18786: data <= 'd0; 18787: data <= 'd0; 18788: data <= 'd0; 18789: data <= 'd0; 18790: data <= 'd0; 18791: data <= 'd0; 18792: data <= 'd0; 18793: data <= 'd2; 18794: data <= 'd1; 18795: data <= 'd3; 18796: data <= 'd6; 18797: data <= 'd6; 18798: data <= 'd6; 18799: data <= 'd6; 18800: data <= 'd6; 18801: data <= 'd6; 18802: data <= 'd6; 18803: data <= 'd3; 18804: data <= 'd1; 18805: data <= 'd2; 18806: data <= 'd0; 18807: data <= 'd0; 18808: data <= 'd0; 18809: data <= 'd0; 18810: data <= 'd0; 18811: data <= 'd0; 18812: data <= 'd0; 18813: data <= 'd0; 18814: data <= 'd0; 18815: data <= 'd0; 18816: data <= 'd0; 18817: data <= 'd0; 18818: data <= 'd0; 18819: data <= 'd0; 18820: data <= 'd0; 18821: data <= 'd0; 18822: data <= 'd0; 18823: data <= 'd0; 18824: data <= 'd0; 18825: data <= 'd2; 18826: data <= 'd1; 18827: data <= 'd3; 18828: data <= 'd3; 18829: data <= 'd6; 18830: data <= 'd6; 18831: data <= 'd6; 18832: data <= 'd6; 18833: data <= 'd6; 18834: data <= 'd3; 18835: data <= 'd3; 18836: data <= 'd1; 18837: data <= 'd2; 18838: data <= 'd0; 18839: data <= 'd0; 18840: data <= 'd0; 18841: data <= 'd0; 18842: data <= 'd0; 18843: data <= 'd0; 18844: data <= 'd0; 18845: data <= 'd0; 18846: data <= 'd0; 18847: data <= 'd0; 18848: data <= 'd0; 18849: data <= 'd0; 18850: data <= 'd0; 18851: data <= 'd0; 18852: data <= 'd0; 18853: data <= 'd0; 18854: data <= 'd0; 18855: data <= 'd0; 18856: data <= 'd2; 18857: data <= 'd1; 18858: data <= 'd1; 18859: data <= 'd1; 18860: data <= 'd3; 18861: data <= 'd3; 18862: data <= 'd3; 18863: data <= 'd3; 18864: data <= 'd3; 18865: data <= 'd3; 18866: data <= 'd3; 18867: data <= 'd1; 18868: data <= 'd1; 18869: data <= 'd1; 18870: data <= 'd2; 18871: data <= 'd0; 18872: data <= 'd0; 18873: data <= 'd0; 18874: data <= 'd0; 18875: data <= 'd0; 18876: data <= 'd0; 18877: data <= 'd0; 18878: data <= 'd0; 18879: data <= 'd0; 18880: data <= 'd0; 18881: data <= 'd0; 18882: data <= 'd0; 18883: data <= 'd0; 18884: data <= 'd0; 18885: data <= 'd0; 18886: data <= 'd0; 18887: data <= 'd0; 18888: data <= 'd5; 18889: data <= 'd5; 18890: data <= 'd1; 18891: data <= 'd3; 18892: data <= 'd3; 18893: data <= 'd3; 18894: data <= 'd3; 18895: data <= 'd3; 18896: data <= 'd3; 18897: data <= 'd3; 18898: data <= 'd3; 18899: data <= 'd3; 18900: data <= 'd1; 18901: data <= 'd5; 18902: data <= 'd5; 18903: data <= 'd0; 18904: data <= 'd0; 18905: data <= 'd0; 18906: data <= 'd0; 18907: data <= 'd0; 18908: data <= 'd0; 18909: data <= 'd0; 18910: data <= 'd0; 18911: data <= 'd0; 18912: data <= 'd0; 18913: data <= 'd0; 18914: data <= 'd0; 18915: data <= 'd0; 18916: data <= 'd0; 18917: data <= 'd0; 18918: data <= 'd0; 18919: data <= 'd2; 18920: data <= 'd3; 18921: data <= 'd3; 18922: data <= 'd1; 18923: data <= 'd3; 18924: data <= 'd3; 18925: data <= 'd3; 18926: data <= 'd3; 18927: data <= 'd6; 18928: data <= 'd3; 18929: data <= 'd3; 18930: data <= 'd3; 18931: data <= 'd3; 18932: data <= 'd1; 18933: data <= 'd3; 18934: data <= 'd3; 18935: data <= 'd2; 18936: data <= 'd0; 18937: data <= 'd0; 18938: data <= 'd0; 18939: data <= 'd0; 18940: data <= 'd0; 18941: data <= 'd0; 18942: data <= 'd0; 18943: data <= 'd0; 18944: data <= 'd0; 18945: data <= 'd0; 18946: data <= 'd0; 18947: data <= 'd0; 18948: data <= 'd0; 18949: data <= 'd0; 18950: data <= 'd0; 18951: data <= 'd2; 18952: data <= 'd3; 18953: data <= 'd3; 18954: data <= 'd3; 18955: data <= 'd1; 18956: data <= 'd3; 18957: data <= 'd3; 18958: data <= 'd6; 18959: data <= 'd6; 18960: data <= 'd6; 18961: data <= 'd3; 18962: data <= 'd3; 18963: data <= 'd1; 18964: data <= 'd3; 18965: data <= 'd3; 18966: data <= 'd3; 18967: data <= 'd2; 18968: data <= 'd0; 18969: data <= 'd0; 18970: data <= 'd0; 18971: data <= 'd0; 18972: data <= 'd0; 18973: data <= 'd0; 18974: data <= 'd0; 18975: data <= 'd0; 18976: data <= 'd0; 18977: data <= 'd0; 18978: data <= 'd0; 18979: data <= 'd0; 18980: data <= 'd0; 18981: data <= 'd0; 18982: data <= 'd0; 18983: data <= 'd2; 18984: data <= 'd1; 18985: data <= 'd1; 18986: data <= 'd3; 18987: data <= 'd1; 18988: data <= 'd5; 18989: data <= 'd3; 18990: data <= 'd6; 18991: data <= 'd6; 18992: data <= 'd6; 18993: data <= 'd3; 18994: data <= 'd5; 18995: data <= 'd1; 18996: data <= 'd3; 18997: data <= 'd1; 18998: data <= 'd1; 18999: data <= 'd2; 19000: data <= 'd0; 19001: data <= 'd0; 19002: data <= 'd0; 19003: data <= 'd0; 19004: data <= 'd0; 19005: data <= 'd0; 19006: data <= 'd0; 19007: data <= 'd0; 19008: data <= 'd0; 19009: data <= 'd0; 19010: data <= 'd0; 19011: data <= 'd0; 19012: data <= 'd0; 19013: data <= 'd0; 19014: data <= 'd0; 19015: data <= 'd0; 19016: data <= 'd2; 19017: data <= 'd2; 19018: data <= 'd1; 19019: data <= 'd1; 19020: data <= 'd5; 19021: data <= 'd3; 19022: data <= 'd3; 19023: data <= 'd6; 19024: data <= 'd3; 19025: data <= 'd3; 19026: data <= 'd5; 19027: data <= 'd1; 19028: data <= 'd1; 19029: data <= 'd2; 19030: data <= 'd2; 19031: data <= 'd0; 19032: data <= 'd0; 19033: data <= 'd0; 19034: data <= 'd0; 19035: data <= 'd0; 19036: data <= 'd0; 19037: data <= 'd0; 19038: data <= 'd0; 19039: data <= 'd0; 19040: data <= 'd0; 19041: data <= 'd0; 19042: data <= 'd0; 19043: data <= 'd0; 19044: data <= 'd0; 19045: data <= 'd0; 19046: data <= 'd0; 19047: data <= 'd0; 19048: data <= 'd2; 19049: data <= 'd8; 19050: data <= 'd2; 19051: data <= 'd2; 19052: data <= 'd2; 19053: data <= 'd1; 19054: data <= 'd3; 19055: data <= 'd3; 19056: data <= 'd3; 19057: data <= 'd1; 19058: data <= 'd2; 19059: data <= 'd2; 19060: data <= 'd2; 19061: data <= 'd8; 19062: data <= 'd2; 19063: data <= 'd0; 19064: data <= 'd0; 19065: data <= 'd0; 19066: data <= 'd0; 19067: data <= 'd0; 19068: data <= 'd0; 19069: data <= 'd0; 19070: data <= 'd0; 19071: data <= 'd0; 19072: data <= 'd0; 19073: data <= 'd0; 19074: data <= 'd0; 19075: data <= 'd0; 19076: data <= 'd0; 19077: data <= 'd0; 19078: data <= 'd0; 19079: data <= 'd0; 19080: data <= 'd0; 19081: data <= 'd2; 19082: data <= 'd8; 19083: data <= 'd8; 19084: data <= 'd2; 19085: data <= 'd1; 19086: data <= 'd3; 19087: data <= 'd3; 19088: data <= 'd3; 19089: data <= 'd1; 19090: data <= 'd2; 19091: data <= 'd8; 19092: data <= 'd8; 19093: data <= 'd2; 19094: data <= 'd0; 19095: data <= 'd0; 19096: data <= 'd0; 19097: data <= 'd0; 19098: data <= 'd0; 19099: data <= 'd0; 19100: data <= 'd0; 19101: data <= 'd0; 19102: data <= 'd0; 19103: data <= 'd0; 19104: data <= 'd0; 19105: data <= 'd0; 19106: data <= 'd0; 19107: data <= 'd0; 19108: data <= 'd0; 19109: data <= 'd0; 19110: data <= 'd0; 19111: data <= 'd0; 19112: data <= 'd0; 19113: data <= 'd2; 19114: data <= 'd9; 19115: data <= 'd8; 19116: data <= 'd8; 19117: data <= 'd2; 19118: data <= 'd1; 19119: data <= 'd3; 19120: data <= 'd1; 19121: data <= 'd2; 19122: data <= 'd8; 19123: data <= 'd8; 19124: data <= 'd9; 19125: data <= 'd2; 19126: data <= 'd0; 19127: data <= 'd0; 19128: data <= 'd0; 19129: data <= 'd0; 19130: data <= 'd0; 19131: data <= 'd0; 19132: data <= 'd0; 19133: data <= 'd0; 19134: data <= 'd0; 19135: data <= 'd0; 19136: data <= 'd0; 19137: data <= 'd0; 19138: data <= 'd0; 19139: data <= 'd0; 19140: data <= 'd0; 19141: data <= 'd0; 19142: data <= 'd0; 19143: data <= 'd0; 19144: data <= 'd0; 19145: data <= 'd2; 19146: data <= 'd2; 19147: data <= 'd8; 19148: data <= 'd8; 19149: data <= 'd8; 19150: data <= 'd2; 19151: data <= 'd2; 19152: data <= 'd2; 19153: data <= 'd8; 19154: data <= 'd8; 19155: data <= 'd9; 19156: data <= 'd8; 19157: data <= 'd2; 19158: data <= 'd0; 19159: data <= 'd0; 19160: data <= 'd0; 19161: data <= 'd0; 19162: data <= 'd0; 19163: data <= 'd0; 19164: data <= 'd0; 19165: data <= 'd0; 19166: data <= 'd0; 19167: data <= 'd0; 19168: data <= 'd0; 19169: data <= 'd0; 19170: data <= 'd0; 19171: data <= 'd0; 19172: data <= 'd0; 19173: data <= 'd0; 19174: data <= 'd0; 19175: data <= 'd0; 19176: data <= 'd2; 19177: data <= 'd4; 19178: data <= 'd7; 19179: data <= 'd1; 19180: data <= 'd3; 19181: data <= 'd3; 19182: data <= 'd1; 19183: data <= 'd1; 19184: data <= 'd1; 19185: data <= 'd3; 19186: data <= 'd3; 19187: data <= 'd1; 19188: data <= 'd7; 19189: data <= 'd4; 19190: data <= 'd2; 19191: data <= 'd0; 19192: data <= 'd0; 19193: data <= 'd0; 19194: data <= 'd0; 19195: data <= 'd0; 19196: data <= 'd0; 19197: data <= 'd0; 19198: data <= 'd0; 19199: data <= 'd0; 19200: data <= 'd0; 19201: data <= 'd0; 19202: data <= 'd0; 19203: data <= 'd0; 19204: data <= 'd0; 19205: data <= 'd0; 19206: data <= 'd0; 19207: data <= 'd0; 19208: data <= 'd2; 19209: data <= 'd9; 19210: data <= 'd7; 19211: data <= 'd5; 19212: data <= 'd3; 19213: data <= 'd3; 19214: data <= 'd3; 19215: data <= 'd3; 19216: data <= 'd3; 19217: data <= 'd3; 19218: data <= 'd3; 19219: data <= 'd5; 19220: data <= 'd7; 19221: data <= 'd9; 19222: data <= 'd2; 19223: data <= 'd0; 19224: data <= 'd0; 19225: data <= 'd0; 19226: data <= 'd0; 19227: data <= 'd0; 19228: data <= 'd0; 19229: data <= 'd0; 19230: data <= 'd0; 19231: data <= 'd0; 19232: data <= 'd0; 19233: data <= 'd0; 19234: data <= 'd0; 19235: data <= 'd0; 19236: data <= 'd0; 19237: data <= 'd0; 19238: data <= 'd0; 19239: data <= 'd0; 19240: data <= 'd2; 19241: data <= 'd9; 19242: data <= 'd4; 19243: data <= 'd1; 19244: data <= 'd3; 19245: data <= 'd3; 19246: data <= 'd3; 19247: data <= 'd3; 19248: data <= 'd3; 19249: data <= 'd3; 19250: data <= 'd3; 19251: data <= 'd1; 19252: data <= 'd4; 19253: data <= 'd9; 19254: data <= 'd2; 19255: data <= 'd0; 19256: data <= 'd0; 19257: data <= 'd0; 19258: data <= 'd0; 19259: data <= 'd0; 19260: data <= 'd0; 19261: data <= 'd0; 19262: data <= 'd0; 19263: data <= 'd0; 19264: data <= 'd0; 19265: data <= 'd0; 19266: data <= 'd0; 19267: data <= 'd0; 19268: data <= 'd0; 19269: data <= 'd0; 19270: data <= 'd0; 19271: data <= 'd0; 19272: data <= 'd0; 19273: data <= 'd2; 19274: data <= 'd2; 19275: data <= 'd1; 19276: data <= 'd1; 19277: data <= 'd3; 19278: data <= 'd3; 19279: data <= 'd3; 19280: data <= 'd3; 19281: data <= 'd3; 19282: data <= 'd1; 19283: data <= 'd1; 19284: data <= 'd2; 19285: data <= 'd2; 19286: data <= 'd0; 19287: data <= 'd0; 19288: data <= 'd0; 19289: data <= 'd0; 19290: data <= 'd0; 19291: data <= 'd0; 19292: data <= 'd0; 19293: data <= 'd0; 19294: data <= 'd0; 19295: data <= 'd0; 19296: data <= 'd0; 19297: data <= 'd0; 19298: data <= 'd0; 19299: data <= 'd0; 19300: data <= 'd0; 19301: data <= 'd0; 19302: data <= 'd0; 19303: data <= 'd0; 19304: data <= 'd0; 19305: data <= 'd0; 19306: data <= 'd2; 19307: data <= 'd2; 19308: data <= 'd2; 19309: data <= 'd2; 19310: data <= 'd5; 19311: data <= 'd5; 19312: data <= 'd5; 19313: data <= 'd2; 19314: data <= 'd2; 19315: data <= 'd2; 19316: data <= 'd2; 19317: data <= 'd0; 19318: data <= 'd0; 19319: data <= 'd0; 19320: data <= 'd0; 19321: data <= 'd0; 19322: data <= 'd0; 19323: data <= 'd0; 19324: data <= 'd0; 19325: data <= 'd0; 19326: data <= 'd0; 19327: data <= 'd0; 19328: data <= 'd0; 19329: data <= 'd0; 19330: data <= 'd0; 19331: data <= 'd0; 19332: data <= 'd0; 19333: data <= 'd0; 19334: data <= 'd0; 19335: data <= 'd0; 19336: data <= 'd0; 19337: data <= 'd0; 19338: data <= 'd2; 19339: data <= 'd1; 19340: data <= 'd1; 19341: data <= 'd3; 19342: data <= 'd3; 19343: data <= 'd3; 19344: data <= 'd3; 19345: data <= 'd3; 19346: data <= 'd1; 19347: data <= 'd1; 19348: data <= 'd2; 19349: data <= 'd0; 19350: data <= 'd0; 19351: data <= 'd0; 19352: data <= 'd0; 19353: data <= 'd0; 19354: data <= 'd0; 19355: data <= 'd0; 19356: data <= 'd0; 19357: data <= 'd0; 19358: data <= 'd0; 19359: data <= 'd0; 19360: data <= 'd0; 19361: data <= 'd0; 19362: data <= 'd0; 19363: data <= 'd0; 19364: data <= 'd0; 19365: data <= 'd0; 19366: data <= 'd0; 19367: data <= 'd0; 19368: data <= 'd0; 19369: data <= 'd0; 19370: data <= 'd2; 19371: data <= 'd7; 19372: data <= 'd7; 19373: data <= 'd4; 19374: data <= 'd2; 19375: data <= 'd2; 19376: data <= 'd2; 19377: data <= 'd4; 19378: data <= 'd7; 19379: data <= 'd7; 19380: data <= 'd2; 19381: data <= 'd0; 19382: data <= 'd0; 19383: data <= 'd0; 19384: data <= 'd0; 19385: data <= 'd0; 19386: data <= 'd0; 19387: data <= 'd0; 19388: data <= 'd0; 19389: data <= 'd0; 19390: data <= 'd0; 19391: data <= 'd0; 19392: data <= 'd0; 19393: data <= 'd0; 19394: data <= 'd0; 19395: data <= 'd0; 19396: data <= 'd0; 19397: data <= 'd0; 19398: data <= 'd0; 19399: data <= 'd0; 19400: data <= 'd0; 19401: data <= 'd0; 19402: data <= 'd2; 19403: data <= 'd7; 19404: data <= 'd4; 19405: data <= 'd2; 19406: data <= 'd0; 19407: data <= 'd0; 19408: data <= 'd0; 19409: data <= 'd2; 19410: data <= 'd4; 19411: data <= 'd7; 19412: data <= 'd2; 19413: data <= 'd0; 19414: data <= 'd0; 19415: data <= 'd0; 19416: data <= 'd0; 19417: data <= 'd0; 19418: data <= 'd0; 19419: data <= 'd0; 19420: data <= 'd0; 19421: data <= 'd0; 19422: data <= 'd0; 19423: data <= 'd0; 19424: data <= 'd0; 19425: data <= 'd0; 19426: data <= 'd0; 19427: data <= 'd0; 19428: data <= 'd0; 19429: data <= 'd0; 19430: data <= 'd0; 19431: data <= 'd0; 19432: data <= 'd0; 19433: data <= 'd0; 19434: data <= 'd2; 19435: data <= 'd2; 19436: data <= 'd2; 19437: data <= 'd0; 19438: data <= 'd0; 19439: data <= 'd0; 19440: data <= 'd0; 19441: data <= 'd0; 19442: data <= 'd2; 19443: data <= 'd2; 19444: data <= 'd2; 19445: data <= 'd0; 19446: data <= 'd0; 19447: data <= 'd0; 19448: data <= 'd0; 19449: data <= 'd0; 19450: data <= 'd0; 19451: data <= 'd0; 19452: data <= 'd0; 19453: data <= 'd0; 19454: data <= 'd0; 19455: data <= 'd0; 19456: data <= 'd0; 19457: data <= 'd0; 19458: data <= 'd0; 19459: data <= 'd0; 19460: data <= 'd0; 19461: data <= 'd0; 19462: data <= 'd0; 19463: data <= 'd0; 19464: data <= 'd0; 19465: data <= 'd0; 19466: data <= 'd0; 19467: data <= 'd0; 19468: data <= 'd0; 19469: data <= 'd0; 19470: data <= 'd0; 19471: data <= 'd0; 19472: data <= 'd0; 19473: data <= 'd0; 19474: data <= 'd0; 19475: data <= 'd0; 19476: data <= 'd0; 19477: data <= 'd0; 19478: data <= 'd0; 19479: data <= 'd0; 19480: data <= 'd0; 19481: data <= 'd0; 19482: data <= 'd0; 19483: data <= 'd0; 19484: data <= 'd0; 19485: data <= 'd0; 19486: data <= 'd0; 19487: data <= 'd0; 19488: data <= 'd0; 19489: data <= 'd0; 19490: data <= 'd0; 19491: data <= 'd0; 19492: data <= 'd0; 19493: data <= 'd0; 19494: data <= 'd0; 19495: data <= 'd0; 19496: data <= 'd0; 19497: data <= 'd0; 19498: data <= 'd0; 19499: data <= 'd0; 19500: data <= 'd0; 19501: data <= 'd0; 19502: data <= 'd0; 19503: data <= 'd0; 19504: data <= 'd0; 19505: data <= 'd0; 19506: data <= 'd0; 19507: data <= 'd0; 19508: data <= 'd0; 19509: data <= 'd0; 19510: data <= 'd0; 19511: data <= 'd0; 19512: data <= 'd0; 19513: data <= 'd0; 19514: data <= 'd0; 19515: data <= 'd0; 19516: data <= 'd0; 19517: data <= 'd0; 19518: data <= 'd0; 19519: data <= 'd0; 19520: data <= 'd0; 19521: data <= 'd0; 19522: data <= 'd0; 19523: data <= 'd0; 19524: data <= 'd0; 19525: data <= 'd0; 19526: data <= 'd0; 19527: data <= 'd0; 19528: data <= 'd0; 19529: data <= 'd0; 19530: data <= 'd0; 19531: data <= 'd0; 19532: data <= 'd0; 19533: data <= 'd0; 19534: data <= 'd0; 19535: data <= 'd0; 19536: data <= 'd0; 19537: data <= 'd0; 19538: data <= 'd0; 19539: data <= 'd0; 19540: data <= 'd0; 19541: data <= 'd0; 19542: data <= 'd0; 19543: data <= 'd0; 19544: data <= 'd0; 19545: data <= 'd0; 19546: data <= 'd0; 19547: data <= 'd0; 19548: data <= 'd0; 19549: data <= 'd0; 19550: data <= 'd0; 19551: data <= 'd0; 19552: data <= 'd0; 19553: data <= 'd0; 19554: data <= 'd0; 19555: data <= 'd0; 19556: data <= 'd0; 19557: data <= 'd0; 19558: data <= 'd0; 19559: data <= 'd0; 19560: data <= 'd0; 19561: data <= 'd0; 19562: data <= 'd0; 19563: data <= 'd0; 19564: data <= 'd0; 19565: data <= 'd0; 19566: data <= 'd0; 19567: data <= 'd0; 19568: data <= 'd0; 19569: data <= 'd0; 19570: data <= 'd0; 19571: data <= 'd0; 19572: data <= 'd0; 19573: data <= 'd0; 19574: data <= 'd0; 19575: data <= 'd0; 19576: data <= 'd0; 19577: data <= 'd0; 19578: data <= 'd0; 19579: data <= 'd0; 19580: data <= 'd0; 19581: data <= 'd0; 19582: data <= 'd0; 19583: data <= 'd0; 19584: data <= 'd0; 19585: data <= 'd0; 19586: data <= 'd0; 19587: data <= 'd0; 19588: data <= 'd0; 19589: data <= 'd0; 19590: data <= 'd0; 19591: data <= 'd0; 19592: data <= 'd0; 19593: data <= 'd0; 19594: data <= 'd0; 19595: data <= 'd0; 19596: data <= 'd0; 19597: data <= 'd0; 19598: data <= 'd0; 19599: data <= 'd0; 19600: data <= 'd0; 19601: data <= 'd0; 19602: data <= 'd0; 19603: data <= 'd0; 19604: data <= 'd0; 19605: data <= 'd0; 19606: data <= 'd0; 19607: data <= 'd0; 19608: data <= 'd0; 19609: data <= 'd0; 19610: data <= 'd0; 19611: data <= 'd0; 19612: data <= 'd0; 19613: data <= 'd0; 19614: data <= 'd0; 19615: data <= 'd0; 19616: data <= 'd0; 19617: data <= 'd0; 19618: data <= 'd0; 19619: data <= 'd0; 19620: data <= 'd0; 19621: data <= 'd0; 19622: data <= 'd0; 19623: data <= 'd0; 19624: data <= 'd0; 19625: data <= 'd0; 19626: data <= 'd0; 19627: data <= 'd0; 19628: data <= 'd0; 19629: data <= 'd0; 19630: data <= 'd0; 19631: data <= 'd0; 19632: data <= 'd0; 19633: data <= 'd0; 19634: data <= 'd0; 19635: data <= 'd0; 19636: data <= 'd0; 19637: data <= 'd0; 19638: data <= 'd0; 19639: data <= 'd0; 19640: data <= 'd0; 19641: data <= 'd0; 19642: data <= 'd0; 19643: data <= 'd0; 19644: data <= 'd0; 19645: data <= 'd0; 19646: data <= 'd0; 19647: data <= 'd0; 19648: data <= 'd0; 19649: data <= 'd0; 19650: data <= 'd0; 19651: data <= 'd0; 19652: data <= 'd0; 19653: data <= 'd0; 19654: data <= 'd0; 19655: data <= 'd0; 19656: data <= 'd0; 19657: data <= 'd0; 19658: data <= 'd0; 19659: data <= 'd0; 19660: data <= 'd0; 19661: data <= 'd0; 19662: data <= 'd0; 19663: data <= 'd0; 19664: data <= 'd0; 19665: data <= 'd0; 19666: data <= 'd0; 19667: data <= 'd0; 19668: data <= 'd0; 19669: data <= 'd0; 19670: data <= 'd0; 19671: data <= 'd0; 19672: data <= 'd0; 19673: data <= 'd0; 19674: data <= 'd0; 19675: data <= 'd0; 19676: data <= 'd0; 19677: data <= 'd0; 19678: data <= 'd0; 19679: data <= 'd0; 19680: data <= 'd0; 19681: data <= 'd0; 19682: data <= 'd0; 19683: data <= 'd0; 19684: data <= 'd0; 19685: data <= 'd0; 19686: data <= 'd0; 19687: data <= 'd0; 19688: data <= 'd0; 19689: data <= 'd0; 19690: data <= 'd0; 19691: data <= 'd0; 19692: data <= 'd0; 19693: data <= 'd0; 19694: data <= 'd0; 19695: data <= 'd0; 19696: data <= 'd0; 19697: data <= 'd0; 19698: data <= 'd0; 19699: data <= 'd0; 19700: data <= 'd0; 19701: data <= 'd0; 19702: data <= 'd0; 19703: data <= 'd0; 19704: data <= 'd0; 19705: data <= 'd0; 19706: data <= 'd0; 19707: data <= 'd0; 19708: data <= 'd0; 19709: data <= 'd0; 19710: data <= 'd0; 19711: data <= 'd0; 19712: data <= 'd0; 19713: data <= 'd0; 19714: data <= 'd0; 19715: data <= 'd0; 19716: data <= 'd0; 19717: data <= 'd0; 19718: data <= 'd0; 19719: data <= 'd0; 19720: data <= 'd0; 19721: data <= 'd0; 19722: data <= 'd0; 19723: data <= 'd0; 19724: data <= 'd0; 19725: data <= 'd2; 19726: data <= 'd2; 19727: data <= 'd2; 19728: data <= 'd2; 19729: data <= 'd2; 19730: data <= 'd0; 19731: data <= 'd0; 19732: data <= 'd0; 19733: data <= 'd0; 19734: data <= 'd0; 19735: data <= 'd0; 19736: data <= 'd0; 19737: data <= 'd0; 19738: data <= 'd0; 19739: data <= 'd0; 19740: data <= 'd0; 19741: data <= 'd0; 19742: data <= 'd0; 19743: data <= 'd0; 19744: data <= 'd0; 19745: data <= 'd0; 19746: data <= 'd0; 19747: data <= 'd0; 19748: data <= 'd0; 19749: data <= 'd0; 19750: data <= 'd0; 19751: data <= 'd0; 19752: data <= 'd0; 19753: data <= 'd0; 19754: data <= 'd0; 19755: data <= 'd2; 19756: data <= 'd2; 19757: data <= 'd6; 19758: data <= 'd6; 19759: data <= 'd6; 19760: data <= 'd6; 19761: data <= 'd6; 19762: data <= 'd2; 19763: data <= 'd2; 19764: data <= 'd0; 19765: data <= 'd0; 19766: data <= 'd0; 19767: data <= 'd0; 19768: data <= 'd0; 19769: data <= 'd0; 19770: data <= 'd0; 19771: data <= 'd0; 19772: data <= 'd0; 19773: data <= 'd0; 19774: data <= 'd0; 19775: data <= 'd0; 19776: data <= 'd0; 19777: data <= 'd0; 19778: data <= 'd0; 19779: data <= 'd0; 19780: data <= 'd0; 19781: data <= 'd0; 19782: data <= 'd0; 19783: data <= 'd0; 19784: data <= 'd0; 19785: data <= 'd0; 19786: data <= 'd2; 19787: data <= 'd3; 19788: data <= 'd6; 19789: data <= 'd6; 19790: data <= 'd6; 19791: data <= 'd6; 19792: data <= 'd6; 19793: data <= 'd6; 19794: data <= 'd6; 19795: data <= 'd3; 19796: data <= 'd2; 19797: data <= 'd0; 19798: data <= 'd0; 19799: data <= 'd0; 19800: data <= 'd0; 19801: data <= 'd0; 19802: data <= 'd0; 19803: data <= 'd0; 19804: data <= 'd0; 19805: data <= 'd0; 19806: data <= 'd0; 19807: data <= 'd0; 19808: data <= 'd0; 19809: data <= 'd0; 19810: data <= 'd0; 19811: data <= 'd0; 19812: data <= 'd0; 19813: data <= 'd0; 19814: data <= 'd0; 19815: data <= 'd0; 19816: data <= 'd0; 19817: data <= 'd2; 19818: data <= 'd1; 19819: data <= 'd3; 19820: data <= 'd6; 19821: data <= 'd6; 19822: data <= 'd6; 19823: data <= 'd6; 19824: data <= 'd6; 19825: data <= 'd6; 19826: data <= 'd6; 19827: data <= 'd3; 19828: data <= 'd1; 19829: data <= 'd2; 19830: data <= 'd0; 19831: data <= 'd0; 19832: data <= 'd0; 19833: data <= 'd0; 19834: data <= 'd0; 19835: data <= 'd0; 19836: data <= 'd0; 19837: data <= 'd0; 19838: data <= 'd0; 19839: data <= 'd0; 19840: data <= 'd0; 19841: data <= 'd0; 19842: data <= 'd0; 19843: data <= 'd0; 19844: data <= 'd0; 19845: data <= 'd0; 19846: data <= 'd0; 19847: data <= 'd0; 19848: data <= 'd0; 19849: data <= 'd2; 19850: data <= 'd1; 19851: data <= 'd3; 19852: data <= 'd3; 19853: data <= 'd6; 19854: data <= 'd6; 19855: data <= 'd6; 19856: data <= 'd6; 19857: data <= 'd6; 19858: data <= 'd3; 19859: data <= 'd3; 19860: data <= 'd1; 19861: data <= 'd2; 19862: data <= 'd0; 19863: data <= 'd0; 19864: data <= 'd0; 19865: data <= 'd0; 19866: data <= 'd0; 19867: data <= 'd0; 19868: data <= 'd0; 19869: data <= 'd0; 19870: data <= 'd0; 19871: data <= 'd0; 19872: data <= 'd0; 19873: data <= 'd0; 19874: data <= 'd0; 19875: data <= 'd0; 19876: data <= 'd0; 19877: data <= 'd0; 19878: data <= 'd0; 19879: data <= 'd0; 19880: data <= 'd2; 19881: data <= 'd1; 19882: data <= 'd1; 19883: data <= 'd1; 19884: data <= 'd3; 19885: data <= 'd3; 19886: data <= 'd3; 19887: data <= 'd3; 19888: data <= 'd3; 19889: data <= 'd3; 19890: data <= 'd3; 19891: data <= 'd1; 19892: data <= 'd1; 19893: data <= 'd1; 19894: data <= 'd2; 19895: data <= 'd0; 19896: data <= 'd0; 19897: data <= 'd0; 19898: data <= 'd0; 19899: data <= 'd0; 19900: data <= 'd0; 19901: data <= 'd0; 19902: data <= 'd0; 19903: data <= 'd0; 19904: data <= 'd0; 19905: data <= 'd0; 19906: data <= 'd0; 19907: data <= 'd0; 19908: data <= 'd0; 19909: data <= 'd0; 19910: data <= 'd0; 19911: data <= 'd0; 19912: data <= 'd5; 19913: data <= 'd5; 19914: data <= 'd1; 19915: data <= 'd3; 19916: data <= 'd3; 19917: data <= 'd3; 19918: data <= 'd3; 19919: data <= 'd3; 19920: data <= 'd3; 19921: data <= 'd3; 19922: data <= 'd3; 19923: data <= 'd3; 19924: data <= 'd1; 19925: data <= 'd5; 19926: data <= 'd5; 19927: data <= 'd0; 19928: data <= 'd0; 19929: data <= 'd0; 19930: data <= 'd0; 19931: data <= 'd0; 19932: data <= 'd0; 19933: data <= 'd0; 19934: data <= 'd0; 19935: data <= 'd0; 19936: data <= 'd0; 19937: data <= 'd0; 19938: data <= 'd0; 19939: data <= 'd0; 19940: data <= 'd0; 19941: data <= 'd0; 19942: data <= 'd0; 19943: data <= 'd2; 19944: data <= 'd3; 19945: data <= 'd3; 19946: data <= 'd1; 19947: data <= 'd3; 19948: data <= 'd3; 19949: data <= 'd3; 19950: data <= 'd3; 19951: data <= 'd6; 19952: data <= 'd3; 19953: data <= 'd3; 19954: data <= 'd3; 19955: data <= 'd3; 19956: data <= 'd1; 19957: data <= 'd3; 19958: data <= 'd3; 19959: data <= 'd2; 19960: data <= 'd0; 19961: data <= 'd0; 19962: data <= 'd0; 19963: data <= 'd0; 19964: data <= 'd0; 19965: data <= 'd0; 19966: data <= 'd0; 19967: data <= 'd0; 19968: data <= 'd0; 19969: data <= 'd0; 19970: data <= 'd0; 19971: data <= 'd0; 19972: data <= 'd0; 19973: data <= 'd0; 19974: data <= 'd0; 19975: data <= 'd2; 19976: data <= 'd3; 19977: data <= 'd3; 19978: data <= 'd3; 19979: data <= 'd1; 19980: data <= 'd3; 19981: data <= 'd3; 19982: data <= 'd6; 19983: data <= 'd6; 19984: data <= 'd6; 19985: data <= 'd3; 19986: data <= 'd3; 19987: data <= 'd1; 19988: data <= 'd3; 19989: data <= 'd3; 19990: data <= 'd3; 19991: data <= 'd2; 19992: data <= 'd0; 19993: data <= 'd0; 19994: data <= 'd0; 19995: data <= 'd0; 19996: data <= 'd0; 19997: data <= 'd0; 19998: data <= 'd0; 19999: data <= 'd0; 20000: data <= 'd0; 20001: data <= 'd0; 20002: data <= 'd0; 20003: data <= 'd0; 20004: data <= 'd0; 20005: data <= 'd0; 20006: data <= 'd0; 20007: data <= 'd2; 20008: data <= 'd1; 20009: data <= 'd1; 20010: data <= 'd3; 20011: data <= 'd1; 20012: data <= 'd5; 20013: data <= 'd3; 20014: data <= 'd6; 20015: data <= 'd6; 20016: data <= 'd6; 20017: data <= 'd3; 20018: data <= 'd5; 20019: data <= 'd1; 20020: data <= 'd3; 20021: data <= 'd1; 20022: data <= 'd1; 20023: data <= 'd2; 20024: data <= 'd0; 20025: data <= 'd0; 20026: data <= 'd0; 20027: data <= 'd0; 20028: data <= 'd0; 20029: data <= 'd0; 20030: data <= 'd0; 20031: data <= 'd0; 20032: data <= 'd0; 20033: data <= 'd0; 20034: data <= 'd0; 20035: data <= 'd0; 20036: data <= 'd0; 20037: data <= 'd0; 20038: data <= 'd0; 20039: data <= 'd0; 20040: data <= 'd2; 20041: data <= 'd2; 20042: data <= 'd1; 20043: data <= 'd1; 20044: data <= 'd5; 20045: data <= 'd3; 20046: data <= 'd3; 20047: data <= 'd6; 20048: data <= 'd3; 20049: data <= 'd3; 20050: data <= 'd5; 20051: data <= 'd1; 20052: data <= 'd1; 20053: data <= 'd2; 20054: data <= 'd2; 20055: data <= 'd0; 20056: data <= 'd0; 20057: data <= 'd0; 20058: data <= 'd0; 20059: data <= 'd0; 20060: data <= 'd0; 20061: data <= 'd0; 20062: data <= 'd0; 20063: data <= 'd0; 20064: data <= 'd0; 20065: data <= 'd0; 20066: data <= 'd0; 20067: data <= 'd0; 20068: data <= 'd0; 20069: data <= 'd0; 20070: data <= 'd0; 20071: data <= 'd0; 20072: data <= 'd2; 20073: data <= 'd8; 20074: data <= 'd2; 20075: data <= 'd2; 20076: data <= 'd2; 20077: data <= 'd1; 20078: data <= 'd3; 20079: data <= 'd3; 20080: data <= 'd3; 20081: data <= 'd1; 20082: data <= 'd2; 20083: data <= 'd2; 20084: data <= 'd2; 20085: data <= 'd8; 20086: data <= 'd2; 20087: data <= 'd0; 20088: data <= 'd0; 20089: data <= 'd0; 20090: data <= 'd0; 20091: data <= 'd0; 20092: data <= 'd0; 20093: data <= 'd0; 20094: data <= 'd0; 20095: data <= 'd0; 20096: data <= 'd0; 20097: data <= 'd0; 20098: data <= 'd0; 20099: data <= 'd0; 20100: data <= 'd0; 20101: data <= 'd0; 20102: data <= 'd0; 20103: data <= 'd0; 20104: data <= 'd0; 20105: data <= 'd2; 20106: data <= 'd8; 20107: data <= 'd8; 20108: data <= 'd2; 20109: data <= 'd1; 20110: data <= 'd3; 20111: data <= 'd3; 20112: data <= 'd3; 20113: data <= 'd2; 20114: data <= 'd8; 20115: data <= 'd8; 20116: data <= 'd8; 20117: data <= 'd2; 20118: data <= 'd0; 20119: data <= 'd0; 20120: data <= 'd0; 20121: data <= 'd0; 20122: data <= 'd0; 20123: data <= 'd0; 20124: data <= 'd0; 20125: data <= 'd0; 20126: data <= 'd0; 20127: data <= 'd0; 20128: data <= 'd0; 20129: data <= 'd0; 20130: data <= 'd0; 20131: data <= 'd0; 20132: data <= 'd0; 20133: data <= 'd0; 20134: data <= 'd0; 20135: data <= 'd0; 20136: data <= 'd0; 20137: data <= 'd2; 20138: data <= 'd9; 20139: data <= 'd8; 20140: data <= 'd2; 20141: data <= 'd1; 20142: data <= 'd3; 20143: data <= 'd1; 20144: data <= 'd2; 20145: data <= 'd8; 20146: data <= 'd9; 20147: data <= 'd8; 20148: data <= 'd5; 20149: data <= 'd9; 20150: data <= 'd2; 20151: data <= 'd0; 20152: data <= 'd0; 20153: data <= 'd0; 20154: data <= 'd0; 20155: data <= 'd0; 20156: data <= 'd0; 20157: data <= 'd0; 20158: data <= 'd0; 20159: data <= 'd0; 20160: data <= 'd0; 20161: data <= 'd0; 20162: data <= 'd0; 20163: data <= 'd0; 20164: data <= 'd0; 20165: data <= 'd0; 20166: data <= 'd0; 20167: data <= 'd0; 20168: data <= 'd0; 20169: data <= 'd2; 20170: data <= 'd2; 20171: data <= 'd8; 20172: data <= 'd8; 20173: data <= 'd2; 20174: data <= 'd2; 20175: data <= 'd2; 20176: data <= 'd8; 20177: data <= 'd9; 20178: data <= 'd9; 20179: data <= 'd9; 20180: data <= 'd4; 20181: data <= 'd9; 20182: data <= 'd2; 20183: data <= 'd0; 20184: data <= 'd0; 20185: data <= 'd0; 20186: data <= 'd0; 20187: data <= 'd0; 20188: data <= 'd0; 20189: data <= 'd0; 20190: data <= 'd0; 20191: data <= 'd0; 20192: data <= 'd0; 20193: data <= 'd0; 20194: data <= 'd0; 20195: data <= 'd0; 20196: data <= 'd0; 20197: data <= 'd0; 20198: data <= 'd0; 20199: data <= 'd0; 20200: data <= 'd0; 20201: data <= 'd2; 20202: data <= 'd7; 20203: data <= 'd1; 20204: data <= 'd3; 20205: data <= 'd1; 20206: data <= 'd1; 20207: data <= 'd1; 20208: data <= 'd3; 20209: data <= 'd3; 20210: data <= 'd3; 20211: data <= 'd1; 20212: data <= 'd7; 20213: data <= 'd2; 20214: data <= 'd0; 20215: data <= 'd0; 20216: data <= 'd0; 20217: data <= 'd0; 20218: data <= 'd0; 20219: data <= 'd0; 20220: data <= 'd0; 20221: data <= 'd0; 20222: data <= 'd0; 20223: data <= 'd0; 20224: data <= 'd0; 20225: data <= 'd0; 20226: data <= 'd0; 20227: data <= 'd0; 20228: data <= 'd0; 20229: data <= 'd0; 20230: data <= 'd0; 20231: data <= 'd0; 20232: data <= 'd2; 20233: data <= 'd4; 20234: data <= 'd7; 20235: data <= 'd5; 20236: data <= 'd3; 20237: data <= 'd3; 20238: data <= 'd3; 20239: data <= 'd3; 20240: data <= 'd3; 20241: data <= 'd3; 20242: data <= 'd3; 20243: data <= 'd5; 20244: data <= 'd7; 20245: data <= 'd2; 20246: data <= 'd0; 20247: data <= 'd0; 20248: data <= 'd0; 20249: data <= 'd0; 20250: data <= 'd0; 20251: data <= 'd0; 20252: data <= 'd0; 20253: data <= 'd0; 20254: data <= 'd0; 20255: data <= 'd0; 20256: data <= 'd0; 20257: data <= 'd0; 20258: data <= 'd0; 20259: data <= 'd0; 20260: data <= 'd0; 20261: data <= 'd0; 20262: data <= 'd0; 20263: data <= 'd0; 20264: data <= 'd2; 20265: data <= 'd9; 20266: data <= 'd4; 20267: data <= 'd1; 20268: data <= 'd3; 20269: data <= 'd3; 20270: data <= 'd3; 20271: data <= 'd3; 20272: data <= 'd3; 20273: data <= 'd3; 20274: data <= 'd3; 20275: data <= 'd1; 20276: data <= 'd2; 20277: data <= 'd0; 20278: data <= 'd0; 20279: data <= 'd0; 20280: data <= 'd0; 20281: data <= 'd0; 20282: data <= 'd0; 20283: data <= 'd0; 20284: data <= 'd0; 20285: data <= 'd0; 20286: data <= 'd0; 20287: data <= 'd0; 20288: data <= 'd0; 20289: data <= 'd0; 20290: data <= 'd0; 20291: data <= 'd0; 20292: data <= 'd0; 20293: data <= 'd0; 20294: data <= 'd0; 20295: data <= 'd0; 20296: data <= 'd2; 20297: data <= 'd9; 20298: data <= 'd2; 20299: data <= 'd1; 20300: data <= 'd1; 20301: data <= 'd3; 20302: data <= 'd3; 20303: data <= 'd3; 20304: data <= 'd3; 20305: data <= 'd3; 20306: data <= 'd1; 20307: data <= 'd1; 20308: data <= 'd2; 20309: data <= 'd0; 20310: data <= 'd0; 20311: data <= 'd0; 20312: data <= 'd0; 20313: data <= 'd0; 20314: data <= 'd0; 20315: data <= 'd0; 20316: data <= 'd0; 20317: data <= 'd0; 20318: data <= 'd0; 20319: data <= 'd0; 20320: data <= 'd0; 20321: data <= 'd0; 20322: data <= 'd0; 20323: data <= 'd0; 20324: data <= 'd0; 20325: data <= 'd0; 20326: data <= 'd0; 20327: data <= 'd0; 20328: data <= 'd0; 20329: data <= 'd2; 20330: data <= 'd2; 20331: data <= 'd2; 20332: data <= 'd2; 20333: data <= 'd2; 20334: data <= 'd5; 20335: data <= 'd5; 20336: data <= 'd5; 20337: data <= 'd2; 20338: data <= 'd2; 20339: data <= 'd2; 20340: data <= 'd2; 20341: data <= 'd0; 20342: data <= 'd0; 20343: data <= 'd0; 20344: data <= 'd0; 20345: data <= 'd0; 20346: data <= 'd0; 20347: data <= 'd0; 20348: data <= 'd0; 20349: data <= 'd0; 20350: data <= 'd0; 20351: data <= 'd0; 20352: data <= 'd0; 20353: data <= 'd0; 20354: data <= 'd0; 20355: data <= 'd0; 20356: data <= 'd0; 20357: data <= 'd0; 20358: data <= 'd0; 20359: data <= 'd0; 20360: data <= 'd0; 20361: data <= 'd0; 20362: data <= 'd2; 20363: data <= 'd1; 20364: data <= 'd1; 20365: data <= 'd3; 20366: data <= 'd3; 20367: data <= 'd3; 20368: data <= 'd3; 20369: data <= 'd3; 20370: data <= 'd1; 20371: data <= 'd1; 20372: data <= 'd2; 20373: data <= 'd0; 20374: data <= 'd0; 20375: data <= 'd0; 20376: data <= 'd0; 20377: data <= 'd0; 20378: data <= 'd0; 20379: data <= 'd0; 20380: data <= 'd0; 20381: data <= 'd0; 20382: data <= 'd0; 20383: data <= 'd0; 20384: data <= 'd0; 20385: data <= 'd0; 20386: data <= 'd0; 20387: data <= 'd0; 20388: data <= 'd0; 20389: data <= 'd0; 20390: data <= 'd0; 20391: data <= 'd0; 20392: data <= 'd0; 20393: data <= 'd0; 20394: data <= 'd2; 20395: data <= 'd7; 20396: data <= 'd7; 20397: data <= 'd2; 20398: data <= 'd2; 20399: data <= 'd2; 20400: data <= 'd2; 20401: data <= 'd4; 20402: data <= 'd7; 20403: data <= 'd7; 20404: data <= 'd2; 20405: data <= 'd0; 20406: data <= 'd0; 20407: data <= 'd0; 20408: data <= 'd0; 20409: data <= 'd0; 20410: data <= 'd0; 20411: data <= 'd0; 20412: data <= 'd0; 20413: data <= 'd0; 20414: data <= 'd0; 20415: data <= 'd0; 20416: data <= 'd0; 20417: data <= 'd0; 20418: data <= 'd0; 20419: data <= 'd0; 20420: data <= 'd0; 20421: data <= 'd0; 20422: data <= 'd0; 20423: data <= 'd0; 20424: data <= 'd0; 20425: data <= 'd0; 20426: data <= 'd2; 20427: data <= 'd2; 20428: data <= 'd2; 20429: data <= 'd0; 20430: data <= 'd0; 20431: data <= 'd0; 20432: data <= 'd0; 20433: data <= 'd2; 20434: data <= 'd7; 20435: data <= 'd4; 20436: data <= 'd2; 20437: data <= 'd0; 20438: data <= 'd0; 20439: data <= 'd0; 20440: data <= 'd0; 20441: data <= 'd0; 20442: data <= 'd0; 20443: data <= 'd0; 20444: data <= 'd0; 20445: data <= 'd0; 20446: data <= 'd0; 20447: data <= 'd0; 20448: data <= 'd0; 20449: data <= 'd0; 20450: data <= 'd0; 20451: data <= 'd0; 20452: data <= 'd0; 20453: data <= 'd0; 20454: data <= 'd0; 20455: data <= 'd0; 20456: data <= 'd0; 20457: data <= 'd0; 20458: data <= 'd0; 20459: data <= 'd0; 20460: data <= 'd0; 20461: data <= 'd0; 20462: data <= 'd0; 20463: data <= 'd0; 20464: data <= 'd0; 20465: data <= 'd2; 20466: data <= 'd2; 20467: data <= 'd2; 20468: data <= 'd0; 20469: data <= 'd0; 20470: data <= 'd0; 20471: data <= 'd0; 20472: data <= 'd0; 20473: data <= 'd0; 20474: data <= 'd0; 20475: data <= 'd0; 20476: data <= 'd0; 20477: data <= 'd0; 20478: data <= 'd0; 20479: data <= 'd0; 20480: data <= 'd0; 20481: data <= 'd0; 20482: data <= 'd0; 20483: data <= 'd0; 20484: data <= 'd0; 20485: data <= 'd0; 20486: data <= 'd0; 20487: data <= 'd0; 20488: data <= 'd0; 20489: data <= 'd0; 20490: data <= 'd0; 20491: data <= 'd0; 20492: data <= 'd0; 20493: data <= 'd0; 20494: data <= 'd0; 20495: data <= 'd0; 20496: data <= 'd0; 20497: data <= 'd0; 20498: data <= 'd0; 20499: data <= 'd0; 20500: data <= 'd0; 20501: data <= 'd0; 20502: data <= 'd0; 20503: data <= 'd0; 20504: data <= 'd0; 20505: data <= 'd0; 20506: data <= 'd0; 20507: data <= 'd0; 20508: data <= 'd0; 20509: data <= 'd0; 20510: data <= 'd0; 20511: data <= 'd0; 20512: data <= 'd0; 20513: data <= 'd0; 20514: data <= 'd0; 20515: data <= 'd0; 20516: data <= 'd0; 20517: data <= 'd0; 20518: data <= 'd0; 20519: data <= 'd0; 20520: data <= 'd0; 20521: data <= 'd0; 20522: data <= 'd0; 20523: data <= 'd0; 20524: data <= 'd0; 20525: data <= 'd0; 20526: data <= 'd0; 20527: data <= 'd0; 20528: data <= 'd0; 20529: data <= 'd0; 20530: data <= 'd0; 20531: data <= 'd0; 20532: data <= 'd0; 20533: data <= 'd0; 20534: data <= 'd0; 20535: data <= 'd0; 20536: data <= 'd0; 20537: data <= 'd0; 20538: data <= 'd0; 20539: data <= 'd0; 20540: data <= 'd0; 20541: data <= 'd0; 20542: data <= 'd0; 20543: data <= 'd0; 20544: data <= 'd0; 20545: data <= 'd0; 20546: data <= 'd0; 20547: data <= 'd0; 20548: data <= 'd0; 20549: data <= 'd0; 20550: data <= 'd0; 20551: data <= 'd0; 20552: data <= 'd0; 20553: data <= 'd0; 20554: data <= 'd0; 20555: data <= 'd0; 20556: data <= 'd0; 20557: data <= 'd0; 20558: data <= 'd0; 20559: data <= 'd0; 20560: data <= 'd0; 20561: data <= 'd0; 20562: data <= 'd0; 20563: data <= 'd0; 20564: data <= 'd0; 20565: data <= 'd0; 20566: data <= 'd0; 20567: data <= 'd0; 20568: data <= 'd0; 20569: data <= 'd0; 20570: data <= 'd0; 20571: data <= 'd0; 20572: data <= 'd0; 20573: data <= 'd0; 20574: data <= 'd0; 20575: data <= 'd0; 20576: data <= 'd0; 20577: data <= 'd0; 20578: data <= 'd0; 20579: data <= 'd0; 20580: data <= 'd0; 20581: data <= 'd0; 20582: data <= 'd0; 20583: data <= 'd0; 20584: data <= 'd0; 20585: data <= 'd0; 20586: data <= 'd0; 20587: data <= 'd0; 20588: data <= 'd0; 20589: data <= 'd0; 20590: data <= 'd0; 20591: data <= 'd0; 20592: data <= 'd0; 20593: data <= 'd0; 20594: data <= 'd0; 20595: data <= 'd0; 20596: data <= 'd0; 20597: data <= 'd0; 20598: data <= 'd0; 20599: data <= 'd0; 20600: data <= 'd0; 20601: data <= 'd0; 20602: data <= 'd0; 20603: data <= 'd0; 20604: data <= 'd0; 20605: data <= 'd0; 20606: data <= 'd0; 20607: data <= 'd0; 20608: data <= 'd0; 20609: data <= 'd0; 20610: data <= 'd0; 20611: data <= 'd0; 20612: data <= 'd0; 20613: data <= 'd0; 20614: data <= 'd0; 20615: data <= 'd0; 20616: data <= 'd0; 20617: data <= 'd0; 20618: data <= 'd0; 20619: data <= 'd0; 20620: data <= 'd0; 20621: data <= 'd0; 20622: data <= 'd0; 20623: data <= 'd0; 20624: data <= 'd0; 20625: data <= 'd0; 20626: data <= 'd0; 20627: data <= 'd0; 20628: data <= 'd0; 20629: data <= 'd0; 20630: data <= 'd0; 20631: data <= 'd0; 20632: data <= 'd0; 20633: data <= 'd0; 20634: data <= 'd0; 20635: data <= 'd0; 20636: data <= 'd0; 20637: data <= 'd0; 20638: data <= 'd0; 20639: data <= 'd0; 20640: data <= 'd0; 20641: data <= 'd0; 20642: data <= 'd0; 20643: data <= 'd0; 20644: data <= 'd0; 20645: data <= 'd0; 20646: data <= 'd0; 20647: data <= 'd0; 20648: data <= 'd0; 20649: data <= 'd0; 20650: data <= 'd0; 20651: data <= 'd0; 20652: data <= 'd0; 20653: data <= 'd0; 20654: data <= 'd0; 20655: data <= 'd0; 20656: data <= 'd0; 20657: data <= 'd0; 20658: data <= 'd0; 20659: data <= 'd0; 20660: data <= 'd0; 20661: data <= 'd0; 20662: data <= 'd0; 20663: data <= 'd0; 20664: data <= 'd0; 20665: data <= 'd0; 20666: data <= 'd0; 20667: data <= 'd0; 20668: data <= 'd0; 20669: data <= 'd0; 20670: data <= 'd0; 20671: data <= 'd0; 20672: data <= 'd0; 20673: data <= 'd0; 20674: data <= 'd0; 20675: data <= 'd0; 20676: data <= 'd0; 20677: data <= 'd0; 20678: data <= 'd0; 20679: data <= 'd0; 20680: data <= 'd0; 20681: data <= 'd0; 20682: data <= 'd0; 20683: data <= 'd0; 20684: data <= 'd0; 20685: data <= 'd0; 20686: data <= 'd0; 20687: data <= 'd0; 20688: data <= 'd0; 20689: data <= 'd0; 20690: data <= 'd0; 20691: data <= 'd0; 20692: data <= 'd0; 20693: data <= 'd0; 20694: data <= 'd0; 20695: data <= 'd0; 20696: data <= 'd0; 20697: data <= 'd0; 20698: data <= 'd0; 20699: data <= 'd0; 20700: data <= 'd0; 20701: data <= 'd0; 20702: data <= 'd0; 20703: data <= 'd0; 20704: data <= 'd0; 20705: data <= 'd0; 20706: data <= 'd0; 20707: data <= 'd0; 20708: data <= 'd0; 20709: data <= 'd0; 20710: data <= 'd0; 20711: data <= 'd0; 20712: data <= 'd0; 20713: data <= 'd0; 20714: data <= 'd0; 20715: data <= 'd0; 20716: data <= 'd0; 20717: data <= 'd0; 20718: data <= 'd0; 20719: data <= 'd0; 20720: data <= 'd0; 20721: data <= 'd0; 20722: data <= 'd0; 20723: data <= 'd0; 20724: data <= 'd0; 20725: data <= 'd0; 20726: data <= 'd0; 20727: data <= 'd0; 20728: data <= 'd0; 20729: data <= 'd0; 20730: data <= 'd0; 20731: data <= 'd0; 20732: data <= 'd0; 20733: data <= 'd0; 20734: data <= 'd0; 20735: data <= 'd0; 20736: data <= 'd0; 20737: data <= 'd0; 20738: data <= 'd0; 20739: data <= 'd0; 20740: data <= 'd0; 20741: data <= 'd0; 20742: data <= 'd0; 20743: data <= 'd0; 20744: data <= 'd0; 20745: data <= 'd0; 20746: data <= 'd0; 20747: data <= 'd0; 20748: data <= 'd0; 20749: data <= 'd2; 20750: data <= 'd2; 20751: data <= 'd2; 20752: data <= 'd2; 20753: data <= 'd2; 20754: data <= 'd0; 20755: data <= 'd0; 20756: data <= 'd0; 20757: data <= 'd0; 20758: data <= 'd0; 20759: data <= 'd0; 20760: data <= 'd0; 20761: data <= 'd0; 20762: data <= 'd0; 20763: data <= 'd0; 20764: data <= 'd0; 20765: data <= 'd0; 20766: data <= 'd0; 20767: data <= 'd0; 20768: data <= 'd0; 20769: data <= 'd0; 20770: data <= 'd0; 20771: data <= 'd0; 20772: data <= 'd0; 20773: data <= 'd0; 20774: data <= 'd0; 20775: data <= 'd0; 20776: data <= 'd0; 20777: data <= 'd0; 20778: data <= 'd0; 20779: data <= 'd2; 20780: data <= 'd2; 20781: data <= 'd6; 20782: data <= 'd6; 20783: data <= 'd6; 20784: data <= 'd6; 20785: data <= 'd6; 20786: data <= 'd2; 20787: data <= 'd2; 20788: data <= 'd0; 20789: data <= 'd0; 20790: data <= 'd0; 20791: data <= 'd0; 20792: data <= 'd0; 20793: data <= 'd0; 20794: data <= 'd0; 20795: data <= 'd0; 20796: data <= 'd0; 20797: data <= 'd0; 20798: data <= 'd0; 20799: data <= 'd0; 20800: data <= 'd0; 20801: data <= 'd0; 20802: data <= 'd0; 20803: data <= 'd0; 20804: data <= 'd0; 20805: data <= 'd0; 20806: data <= 'd0; 20807: data <= 'd0; 20808: data <= 'd0; 20809: data <= 'd0; 20810: data <= 'd2; 20811: data <= 'd3; 20812: data <= 'd6; 20813: data <= 'd6; 20814: data <= 'd6; 20815: data <= 'd6; 20816: data <= 'd6; 20817: data <= 'd6; 20818: data <= 'd6; 20819: data <= 'd3; 20820: data <= 'd2; 20821: data <= 'd0; 20822: data <= 'd0; 20823: data <= 'd0; 20824: data <= 'd0; 20825: data <= 'd0; 20826: data <= 'd0; 20827: data <= 'd0; 20828: data <= 'd0; 20829: data <= 'd0; 20830: data <= 'd0; 20831: data <= 'd0; 20832: data <= 'd0; 20833: data <= 'd0; 20834: data <= 'd0; 20835: data <= 'd0; 20836: data <= 'd0; 20837: data <= 'd0; 20838: data <= 'd0; 20839: data <= 'd0; 20840: data <= 'd0; 20841: data <= 'd2; 20842: data <= 'd1; 20843: data <= 'd3; 20844: data <= 'd6; 20845: data <= 'd6; 20846: data <= 'd6; 20847: data <= 'd6; 20848: data <= 'd6; 20849: data <= 'd6; 20850: data <= 'd6; 20851: data <= 'd3; 20852: data <= 'd1; 20853: data <= 'd2; 20854: data <= 'd0; 20855: data <= 'd0; 20856: data <= 'd0; 20857: data <= 'd0; 20858: data <= 'd0; 20859: data <= 'd0; 20860: data <= 'd0; 20861: data <= 'd0; 20862: data <= 'd0; 20863: data <= 'd0; 20864: data <= 'd0; 20865: data <= 'd0; 20866: data <= 'd0; 20867: data <= 'd0; 20868: data <= 'd0; 20869: data <= 'd0; 20870: data <= 'd0; 20871: data <= 'd0; 20872: data <= 'd0; 20873: data <= 'd2; 20874: data <= 'd1; 20875: data <= 'd3; 20876: data <= 'd3; 20877: data <= 'd6; 20878: data <= 'd6; 20879: data <= 'd6; 20880: data <= 'd6; 20881: data <= 'd6; 20882: data <= 'd3; 20883: data <= 'd3; 20884: data <= 'd1; 20885: data <= 'd2; 20886: data <= 'd0; 20887: data <= 'd0; 20888: data <= 'd0; 20889: data <= 'd0; 20890: data <= 'd0; 20891: data <= 'd0; 20892: data <= 'd0; 20893: data <= 'd0; 20894: data <= 'd0; 20895: data <= 'd0; 20896: data <= 'd0; 20897: data <= 'd0; 20898: data <= 'd0; 20899: data <= 'd0; 20900: data <= 'd0; 20901: data <= 'd0; 20902: data <= 'd0; 20903: data <= 'd0; 20904: data <= 'd2; 20905: data <= 'd1; 20906: data <= 'd1; 20907: data <= 'd1; 20908: data <= 'd3; 20909: data <= 'd3; 20910: data <= 'd3; 20911: data <= 'd3; 20912: data <= 'd3; 20913: data <= 'd3; 20914: data <= 'd3; 20915: data <= 'd1; 20916: data <= 'd1; 20917: data <= 'd1; 20918: data <= 'd2; 20919: data <= 'd0; 20920: data <= 'd0; 20921: data <= 'd0; 20922: data <= 'd0; 20923: data <= 'd0; 20924: data <= 'd0; 20925: data <= 'd0; 20926: data <= 'd0; 20927: data <= 'd0; 20928: data <= 'd0; 20929: data <= 'd0; 20930: data <= 'd0; 20931: data <= 'd0; 20932: data <= 'd0; 20933: data <= 'd0; 20934: data <= 'd0; 20935: data <= 'd0; 20936: data <= 'd5; 20937: data <= 'd5; 20938: data <= 'd1; 20939: data <= 'd3; 20940: data <= 'd3; 20941: data <= 'd3; 20942: data <= 'd3; 20943: data <= 'd3; 20944: data <= 'd3; 20945: data <= 'd3; 20946: data <= 'd3; 20947: data <= 'd3; 20948: data <= 'd1; 20949: data <= 'd5; 20950: data <= 'd5; 20951: data <= 'd0; 20952: data <= 'd0; 20953: data <= 'd0; 20954: data <= 'd0; 20955: data <= 'd0; 20956: data <= 'd0; 20957: data <= 'd0; 20958: data <= 'd0; 20959: data <= 'd0; 20960: data <= 'd0; 20961: data <= 'd0; 20962: data <= 'd0; 20963: data <= 'd0; 20964: data <= 'd0; 20965: data <= 'd0; 20966: data <= 'd0; 20967: data <= 'd2; 20968: data <= 'd3; 20969: data <= 'd3; 20970: data <= 'd1; 20971: data <= 'd3; 20972: data <= 'd3; 20973: data <= 'd3; 20974: data <= 'd3; 20975: data <= 'd6; 20976: data <= 'd3; 20977: data <= 'd3; 20978: data <= 'd3; 20979: data <= 'd3; 20980: data <= 'd1; 20981: data <= 'd3; 20982: data <= 'd3; 20983: data <= 'd2; 20984: data <= 'd0; 20985: data <= 'd0; 20986: data <= 'd0; 20987: data <= 'd0; 20988: data <= 'd0; 20989: data <= 'd0; 20990: data <= 'd0; 20991: data <= 'd0; 20992: data <= 'd0; 20993: data <= 'd0; 20994: data <= 'd0; 20995: data <= 'd0; 20996: data <= 'd0; 20997: data <= 'd0; 20998: data <= 'd0; 20999: data <= 'd2; 21000: data <= 'd3; 21001: data <= 'd3; 21002: data <= 'd3; 21003: data <= 'd1; 21004: data <= 'd3; 21005: data <= 'd3; 21006: data <= 'd6; 21007: data <= 'd6; 21008: data <= 'd6; 21009: data <= 'd3; 21010: data <= 'd3; 21011: data <= 'd1; 21012: data <= 'd3; 21013: data <= 'd3; 21014: data <= 'd3; 21015: data <= 'd2; 21016: data <= 'd0; 21017: data <= 'd0; 21018: data <= 'd0; 21019: data <= 'd0; 21020: data <= 'd0; 21021: data <= 'd0; 21022: data <= 'd0; 21023: data <= 'd0; 21024: data <= 'd0; 21025: data <= 'd0; 21026: data <= 'd0; 21027: data <= 'd0; 21028: data <= 'd0; 21029: data <= 'd0; 21030: data <= 'd0; 21031: data <= 'd2; 21032: data <= 'd1; 21033: data <= 'd1; 21034: data <= 'd3; 21035: data <= 'd1; 21036: data <= 'd5; 21037: data <= 'd3; 21038: data <= 'd6; 21039: data <= 'd6; 21040: data <= 'd6; 21041: data <= 'd3; 21042: data <= 'd5; 21043: data <= 'd1; 21044: data <= 'd3; 21045: data <= 'd1; 21046: data <= 'd1; 21047: data <= 'd2; 21048: data <= 'd0; 21049: data <= 'd0; 21050: data <= 'd0; 21051: data <= 'd0; 21052: data <= 'd0; 21053: data <= 'd0; 21054: data <= 'd0; 21055: data <= 'd0; 21056: data <= 'd0; 21057: data <= 'd0; 21058: data <= 'd0; 21059: data <= 'd0; 21060: data <= 'd0; 21061: data <= 'd0; 21062: data <= 'd0; 21063: data <= 'd0; 21064: data <= 'd2; 21065: data <= 'd2; 21066: data <= 'd1; 21067: data <= 'd1; 21068: data <= 'd5; 21069: data <= 'd3; 21070: data <= 'd3; 21071: data <= 'd6; 21072: data <= 'd3; 21073: data <= 'd3; 21074: data <= 'd5; 21075: data <= 'd1; 21076: data <= 'd1; 21077: data <= 'd2; 21078: data <= 'd2; 21079: data <= 'd0; 21080: data <= 'd0; 21081: data <= 'd0; 21082: data <= 'd0; 21083: data <= 'd0; 21084: data <= 'd0; 21085: data <= 'd0; 21086: data <= 'd0; 21087: data <= 'd0; 21088: data <= 'd0; 21089: data <= 'd0; 21090: data <= 'd0; 21091: data <= 'd0; 21092: data <= 'd0; 21093: data <= 'd0; 21094: data <= 'd0; 21095: data <= 'd0; 21096: data <= 'd2; 21097: data <= 'd8; 21098: data <= 'd2; 21099: data <= 'd2; 21100: data <= 'd2; 21101: data <= 'd1; 21102: data <= 'd3; 21103: data <= 'd3; 21104: data <= 'd3; 21105: data <= 'd1; 21106: data <= 'd2; 21107: data <= 'd2; 21108: data <= 'd2; 21109: data <= 'd8; 21110: data <= 'd2; 21111: data <= 'd0; 21112: data <= 'd0; 21113: data <= 'd0; 21114: data <= 'd0; 21115: data <= 'd0; 21116: data <= 'd0; 21117: data <= 'd0; 21118: data <= 'd0; 21119: data <= 'd0; 21120: data <= 'd0; 21121: data <= 'd0; 21122: data <= 'd0; 21123: data <= 'd0; 21124: data <= 'd0; 21125: data <= 'd0; 21126: data <= 'd0; 21127: data <= 'd0; 21128: data <= 'd0; 21129: data <= 'd2; 21130: data <= 'd8; 21131: data <= 'd8; 21132: data <= 'd2; 21133: data <= 'd1; 21134: data <= 'd3; 21135: data <= 'd3; 21136: data <= 'd3; 21137: data <= 'd1; 21138: data <= 'd2; 21139: data <= 'd8; 21140: data <= 'd8; 21141: data <= 'd2; 21142: data <= 'd0; 21143: data <= 'd0; 21144: data <= 'd0; 21145: data <= 'd0; 21146: data <= 'd0; 21147: data <= 'd0; 21148: data <= 'd0; 21149: data <= 'd0; 21150: data <= 'd0; 21151: data <= 'd0; 21152: data <= 'd0; 21153: data <= 'd0; 21154: data <= 'd0; 21155: data <= 'd0; 21156: data <= 'd0; 21157: data <= 'd0; 21158: data <= 'd0; 21159: data <= 'd0; 21160: data <= 'd0; 21161: data <= 'd2; 21162: data <= 'd9; 21163: data <= 'd8; 21164: data <= 'd8; 21165: data <= 'd2; 21166: data <= 'd1; 21167: data <= 'd3; 21168: data <= 'd1; 21169: data <= 'd2; 21170: data <= 'd8; 21171: data <= 'd8; 21172: data <= 'd9; 21173: data <= 'd2; 21174: data <= 'd0; 21175: data <= 'd0; 21176: data <= 'd0; 21177: data <= 'd0; 21178: data <= 'd0; 21179: data <= 'd0; 21180: data <= 'd0; 21181: data <= 'd0; 21182: data <= 'd0; 21183: data <= 'd0; 21184: data <= 'd0; 21185: data <= 'd0; 21186: data <= 'd0; 21187: data <= 'd0; 21188: data <= 'd0; 21189: data <= 'd0; 21190: data <= 'd0; 21191: data <= 'd0; 21192: data <= 'd0; 21193: data <= 'd2; 21194: data <= 'd2; 21195: data <= 'd8; 21196: data <= 'd8; 21197: data <= 'd8; 21198: data <= 'd2; 21199: data <= 'd2; 21200: data <= 'd2; 21201: data <= 'd8; 21202: data <= 'd8; 21203: data <= 'd9; 21204: data <= 'd8; 21205: data <= 'd2; 21206: data <= 'd0; 21207: data <= 'd0; 21208: data <= 'd0; 21209: data <= 'd0; 21210: data <= 'd0; 21211: data <= 'd0; 21212: data <= 'd0; 21213: data <= 'd0; 21214: data <= 'd0; 21215: data <= 'd0; 21216: data <= 'd0; 21217: data <= 'd0; 21218: data <= 'd0; 21219: data <= 'd0; 21220: data <= 'd0; 21221: data <= 'd0; 21222: data <= 'd0; 21223: data <= 'd0; 21224: data <= 'd2; 21225: data <= 'd4; 21226: data <= 'd7; 21227: data <= 'd1; 21228: data <= 'd3; 21229: data <= 'd3; 21230: data <= 'd1; 21231: data <= 'd1; 21232: data <= 'd1; 21233: data <= 'd3; 21234: data <= 'd3; 21235: data <= 'd1; 21236: data <= 'd7; 21237: data <= 'd4; 21238: data <= 'd2; 21239: data <= 'd0; 21240: data <= 'd0; 21241: data <= 'd0; 21242: data <= 'd0; 21243: data <= 'd0; 21244: data <= 'd0; 21245: data <= 'd0; 21246: data <= 'd0; 21247: data <= 'd0; 21248: data <= 'd0; 21249: data <= 'd0; 21250: data <= 'd0; 21251: data <= 'd0; 21252: data <= 'd0; 21253: data <= 'd0; 21254: data <= 'd0; 21255: data <= 'd0; 21256: data <= 'd2; 21257: data <= 'd9; 21258: data <= 'd7; 21259: data <= 'd5; 21260: data <= 'd3; 21261: data <= 'd3; 21262: data <= 'd3; 21263: data <= 'd3; 21264: data <= 'd3; 21265: data <= 'd3; 21266: data <= 'd3; 21267: data <= 'd5; 21268: data <= 'd7; 21269: data <= 'd9; 21270: data <= 'd2; 21271: data <= 'd0; 21272: data <= 'd0; 21273: data <= 'd0; 21274: data <= 'd0; 21275: data <= 'd0; 21276: data <= 'd0; 21277: data <= 'd0; 21278: data <= 'd0; 21279: data <= 'd0; 21280: data <= 'd0; 21281: data <= 'd0; 21282: data <= 'd0; 21283: data <= 'd0; 21284: data <= 'd0; 21285: data <= 'd0; 21286: data <= 'd0; 21287: data <= 'd0; 21288: data <= 'd2; 21289: data <= 'd9; 21290: data <= 'd4; 21291: data <= 'd1; 21292: data <= 'd3; 21293: data <= 'd3; 21294: data <= 'd3; 21295: data <= 'd3; 21296: data <= 'd3; 21297: data <= 'd3; 21298: data <= 'd3; 21299: data <= 'd1; 21300: data <= 'd4; 21301: data <= 'd9; 21302: data <= 'd2; 21303: data <= 'd0; 21304: data <= 'd0; 21305: data <= 'd0; 21306: data <= 'd0; 21307: data <= 'd0; 21308: data <= 'd0; 21309: data <= 'd0; 21310: data <= 'd0; 21311: data <= 'd0; 21312: data <= 'd0; 21313: data <= 'd0; 21314: data <= 'd0; 21315: data <= 'd0; 21316: data <= 'd0; 21317: data <= 'd0; 21318: data <= 'd0; 21319: data <= 'd0; 21320: data <= 'd0; 21321: data <= 'd2; 21322: data <= 'd2; 21323: data <= 'd1; 21324: data <= 'd1; 21325: data <= 'd3; 21326: data <= 'd3; 21327: data <= 'd3; 21328: data <= 'd3; 21329: data <= 'd3; 21330: data <= 'd1; 21331: data <= 'd1; 21332: data <= 'd2; 21333: data <= 'd2; 21334: data <= 'd0; 21335: data <= 'd0; 21336: data <= 'd0; 21337: data <= 'd0; 21338: data <= 'd0; 21339: data <= 'd0; 21340: data <= 'd0; 21341: data <= 'd0; 21342: data <= 'd0; 21343: data <= 'd0; 21344: data <= 'd0; 21345: data <= 'd0; 21346: data <= 'd0; 21347: data <= 'd0; 21348: data <= 'd0; 21349: data <= 'd0; 21350: data <= 'd0; 21351: data <= 'd0; 21352: data <= 'd0; 21353: data <= 'd0; 21354: data <= 'd2; 21355: data <= 'd2; 21356: data <= 'd2; 21357: data <= 'd2; 21358: data <= 'd5; 21359: data <= 'd5; 21360: data <= 'd5; 21361: data <= 'd2; 21362: data <= 'd2; 21363: data <= 'd2; 21364: data <= 'd2; 21365: data <= 'd0; 21366: data <= 'd0; 21367: data <= 'd0; 21368: data <= 'd0; 21369: data <= 'd0; 21370: data <= 'd0; 21371: data <= 'd0; 21372: data <= 'd0; 21373: data <= 'd0; 21374: data <= 'd0; 21375: data <= 'd0; 21376: data <= 'd0; 21377: data <= 'd0; 21378: data <= 'd0; 21379: data <= 'd0; 21380: data <= 'd0; 21381: data <= 'd0; 21382: data <= 'd0; 21383: data <= 'd0; 21384: data <= 'd0; 21385: data <= 'd0; 21386: data <= 'd2; 21387: data <= 'd1; 21388: data <= 'd1; 21389: data <= 'd3; 21390: data <= 'd3; 21391: data <= 'd3; 21392: data <= 'd3; 21393: data <= 'd3; 21394: data <= 'd1; 21395: data <= 'd1; 21396: data <= 'd2; 21397: data <= 'd0; 21398: data <= 'd0; 21399: data <= 'd0; 21400: data <= 'd0; 21401: data <= 'd0; 21402: data <= 'd0; 21403: data <= 'd0; 21404: data <= 'd0; 21405: data <= 'd0; 21406: data <= 'd0; 21407: data <= 'd0; 21408: data <= 'd0; 21409: data <= 'd0; 21410: data <= 'd0; 21411: data <= 'd0; 21412: data <= 'd0; 21413: data <= 'd0; 21414: data <= 'd0; 21415: data <= 'd0; 21416: data <= 'd0; 21417: data <= 'd0; 21418: data <= 'd2; 21419: data <= 'd7; 21420: data <= 'd7; 21421: data <= 'd4; 21422: data <= 'd2; 21423: data <= 'd2; 21424: data <= 'd2; 21425: data <= 'd4; 21426: data <= 'd7; 21427: data <= 'd7; 21428: data <= 'd2; 21429: data <= 'd0; 21430: data <= 'd0; 21431: data <= 'd0; 21432: data <= 'd0; 21433: data <= 'd0; 21434: data <= 'd0; 21435: data <= 'd0; 21436: data <= 'd0; 21437: data <= 'd0; 21438: data <= 'd0; 21439: data <= 'd0; 21440: data <= 'd0; 21441: data <= 'd0; 21442: data <= 'd0; 21443: data <= 'd0; 21444: data <= 'd0; 21445: data <= 'd0; 21446: data <= 'd0; 21447: data <= 'd0; 21448: data <= 'd0; 21449: data <= 'd0; 21450: data <= 'd2; 21451: data <= 'd7; 21452: data <= 'd4; 21453: data <= 'd2; 21454: data <= 'd0; 21455: data <= 'd0; 21456: data <= 'd0; 21457: data <= 'd2; 21458: data <= 'd4; 21459: data <= 'd7; 21460: data <= 'd2; 21461: data <= 'd0; 21462: data <= 'd0; 21463: data <= 'd0; 21464: data <= 'd0; 21465: data <= 'd0; 21466: data <= 'd0; 21467: data <= 'd0; 21468: data <= 'd0; 21469: data <= 'd0; 21470: data <= 'd0; 21471: data <= 'd0; 21472: data <= 'd0; 21473: data <= 'd0; 21474: data <= 'd0; 21475: data <= 'd0; 21476: data <= 'd0; 21477: data <= 'd0; 21478: data <= 'd0; 21479: data <= 'd0; 21480: data <= 'd0; 21481: data <= 'd0; 21482: data <= 'd2; 21483: data <= 'd2; 21484: data <= 'd2; 21485: data <= 'd0; 21486: data <= 'd0; 21487: data <= 'd0; 21488: data <= 'd0; 21489: data <= 'd0; 21490: data <= 'd2; 21491: data <= 'd2; 21492: data <= 'd2; 21493: data <= 'd0; 21494: data <= 'd0; 21495: data <= 'd0; 21496: data <= 'd0; 21497: data <= 'd0; 21498: data <= 'd0; 21499: data <= 'd0; 21500: data <= 'd0; 21501: data <= 'd0; 21502: data <= 'd0; 21503: data <= 'd0; 21504: data <= 'd0; 21505: data <= 'd0; 21506: data <= 'd0; 21507: data <= 'd0; 21508: data <= 'd0; 21509: data <= 'd0; 21510: data <= 'd0; 21511: data <= 'd0; 21512: data <= 'd0; 21513: data <= 'd0; 21514: data <= 'd0; 21515: data <= 'd0; 21516: data <= 'd0; 21517: data <= 'd0; 21518: data <= 'd0; 21519: data <= 'd0; 21520: data <= 'd0; 21521: data <= 'd0; 21522: data <= 'd0; 21523: data <= 'd0; 21524: data <= 'd0; 21525: data <= 'd0; 21526: data <= 'd0; 21527: data <= 'd0; 21528: data <= 'd0; 21529: data <= 'd0; 21530: data <= 'd0; 21531: data <= 'd0; 21532: data <= 'd0; 21533: data <= 'd0; 21534: data <= 'd0; 21535: data <= 'd0; 21536: data <= 'd0; 21537: data <= 'd0; 21538: data <= 'd0; 21539: data <= 'd0; 21540: data <= 'd0; 21541: data <= 'd0; 21542: data <= 'd0; 21543: data <= 'd0; 21544: data <= 'd0; 21545: data <= 'd0; 21546: data <= 'd0; 21547: data <= 'd0; 21548: data <= 'd0; 21549: data <= 'd0; 21550: data <= 'd0; 21551: data <= 'd0; 21552: data <= 'd0; 21553: data <= 'd0; 21554: data <= 'd0; 21555: data <= 'd0; 21556: data <= 'd0; 21557: data <= 'd0; 21558: data <= 'd0; 21559: data <= 'd0; 21560: data <= 'd0; 21561: data <= 'd0; 21562: data <= 'd0; 21563: data <= 'd0; 21564: data <= 'd0; 21565: data <= 'd0; 21566: data <= 'd0; 21567: data <= 'd0; 21568: data <= 'd0; 21569: data <= 'd0; 21570: data <= 'd0; 21571: data <= 'd0; 21572: data <= 'd0; 21573: data <= 'd0; 21574: data <= 'd0; 21575: data <= 'd0; 21576: data <= 'd0; 21577: data <= 'd0; 21578: data <= 'd0; 21579: data <= 'd0; 21580: data <= 'd0; 21581: data <= 'd0; 21582: data <= 'd0; 21583: data <= 'd0; 21584: data <= 'd0; 21585: data <= 'd0; 21586: data <= 'd0; 21587: data <= 'd0; 21588: data <= 'd0; 21589: data <= 'd0; 21590: data <= 'd0; 21591: data <= 'd0; 21592: data <= 'd0; 21593: data <= 'd0; 21594: data <= 'd0; 21595: data <= 'd0; 21596: data <= 'd0; 21597: data <= 'd0; 21598: data <= 'd0; 21599: data <= 'd0; 21600: data <= 'd0; 21601: data <= 'd0; 21602: data <= 'd0; 21603: data <= 'd0; 21604: data <= 'd0; 21605: data <= 'd0; 21606: data <= 'd0; 21607: data <= 'd0; 21608: data <= 'd0; 21609: data <= 'd0; 21610: data <= 'd0; 21611: data <= 'd0; 21612: data <= 'd0; 21613: data <= 'd0; 21614: data <= 'd0; 21615: data <= 'd0; 21616: data <= 'd0; 21617: data <= 'd0; 21618: data <= 'd0; 21619: data <= 'd0; 21620: data <= 'd0; 21621: data <= 'd0; 21622: data <= 'd0; 21623: data <= 'd0; 21624: data <= 'd0; 21625: data <= 'd0; 21626: data <= 'd0; 21627: data <= 'd0; 21628: data <= 'd0; 21629: data <= 'd0; 21630: data <= 'd0; 21631: data <= 'd0; 21632: data <= 'd0; 21633: data <= 'd0; 21634: data <= 'd0; 21635: data <= 'd0; 21636: data <= 'd0; 21637: data <= 'd0; 21638: data <= 'd0; 21639: data <= 'd0; 21640: data <= 'd0; 21641: data <= 'd0; 21642: data <= 'd0; 21643: data <= 'd0; 21644: data <= 'd0; 21645: data <= 'd0; 21646: data <= 'd0; 21647: data <= 'd0; 21648: data <= 'd0; 21649: data <= 'd0; 21650: data <= 'd0; 21651: data <= 'd0; 21652: data <= 'd0; 21653: data <= 'd0; 21654: data <= 'd0; 21655: data <= 'd0; 21656: data <= 'd0; 21657: data <= 'd0; 21658: data <= 'd0; 21659: data <= 'd0; 21660: data <= 'd0; 21661: data <= 'd0; 21662: data <= 'd0; 21663: data <= 'd0; 21664: data <= 'd0; 21665: data <= 'd0; 21666: data <= 'd0; 21667: data <= 'd0; 21668: data <= 'd0; 21669: data <= 'd0; 21670: data <= 'd0; 21671: data <= 'd0; 21672: data <= 'd0; 21673: data <= 'd0; 21674: data <= 'd0; 21675: data <= 'd0; 21676: data <= 'd0; 21677: data <= 'd0; 21678: data <= 'd0; 21679: data <= 'd0; 21680: data <= 'd0; 21681: data <= 'd0; 21682: data <= 'd0; 21683: data <= 'd0; 21684: data <= 'd0; 21685: data <= 'd0; 21686: data <= 'd0; 21687: data <= 'd0; 21688: data <= 'd0; 21689: data <= 'd0; 21690: data <= 'd0; 21691: data <= 'd0; 21692: data <= 'd0; 21693: data <= 'd0; 21694: data <= 'd0; 21695: data <= 'd0; 21696: data <= 'd0; 21697: data <= 'd0; 21698: data <= 'd0; 21699: data <= 'd0; 21700: data <= 'd0; 21701: data <= 'd0; 21702: data <= 'd0; 21703: data <= 'd0; 21704: data <= 'd0; 21705: data <= 'd0; 21706: data <= 'd0; 21707: data <= 'd0; 21708: data <= 'd0; 21709: data <= 'd0; 21710: data <= 'd0; 21711: data <= 'd0; 21712: data <= 'd0; 21713: data <= 'd0; 21714: data <= 'd0; 21715: data <= 'd0; 21716: data <= 'd0; 21717: data <= 'd0; 21718: data <= 'd0; 21719: data <= 'd0; 21720: data <= 'd0; 21721: data <= 'd0; 21722: data <= 'd0; 21723: data <= 'd0; 21724: data <= 'd0; 21725: data <= 'd0; 21726: data <= 'd0; 21727: data <= 'd0; 21728: data <= 'd0; 21729: data <= 'd0; 21730: data <= 'd0; 21731: data <= 'd0; 21732: data <= 'd0; 21733: data <= 'd0; 21734: data <= 'd0; 21735: data <= 'd0; 21736: data <= 'd0; 21737: data <= 'd0; 21738: data <= 'd0; 21739: data <= 'd0; 21740: data <= 'd0; 21741: data <= 'd0; 21742: data <= 'd0; 21743: data <= 'd0; 21744: data <= 'd0; 21745: data <= 'd0; 21746: data <= 'd0; 21747: data <= 'd0; 21748: data <= 'd0; 21749: data <= 'd0; 21750: data <= 'd0; 21751: data <= 'd0; 21752: data <= 'd0; 21753: data <= 'd0; 21754: data <= 'd0; 21755: data <= 'd0; 21756: data <= 'd0; 21757: data <= 'd0; 21758: data <= 'd0; 21759: data <= 'd0; 21760: data <= 'd0; 21761: data <= 'd0; 21762: data <= 'd0; 21763: data <= 'd0; 21764: data <= 'd0; 21765: data <= 'd0; 21766: data <= 'd0; 21767: data <= 'd0; 21768: data <= 'd0; 21769: data <= 'd0; 21770: data <= 'd0; 21771: data <= 'd0; 21772: data <= 'd0; 21773: data <= 'd2; 21774: data <= 'd2; 21775: data <= 'd2; 21776: data <= 'd2; 21777: data <= 'd2; 21778: data <= 'd0; 21779: data <= 'd0; 21780: data <= 'd0; 21781: data <= 'd0; 21782: data <= 'd0; 21783: data <= 'd0; 21784: data <= 'd0; 21785: data <= 'd0; 21786: data <= 'd0; 21787: data <= 'd0; 21788: data <= 'd0; 21789: data <= 'd0; 21790: data <= 'd0; 21791: data <= 'd0; 21792: data <= 'd0; 21793: data <= 'd0; 21794: data <= 'd0; 21795: data <= 'd0; 21796: data <= 'd0; 21797: data <= 'd0; 21798: data <= 'd0; 21799: data <= 'd0; 21800: data <= 'd0; 21801: data <= 'd0; 21802: data <= 'd0; 21803: data <= 'd2; 21804: data <= 'd2; 21805: data <= 'd6; 21806: data <= 'd6; 21807: data <= 'd6; 21808: data <= 'd6; 21809: data <= 'd6; 21810: data <= 'd2; 21811: data <= 'd2; 21812: data <= 'd0; 21813: data <= 'd0; 21814: data <= 'd0; 21815: data <= 'd0; 21816: data <= 'd0; 21817: data <= 'd0; 21818: data <= 'd0; 21819: data <= 'd0; 21820: data <= 'd0; 21821: data <= 'd0; 21822: data <= 'd0; 21823: data <= 'd0; 21824: data <= 'd0; 21825: data <= 'd0; 21826: data <= 'd0; 21827: data <= 'd0; 21828: data <= 'd0; 21829: data <= 'd0; 21830: data <= 'd0; 21831: data <= 'd0; 21832: data <= 'd0; 21833: data <= 'd0; 21834: data <= 'd2; 21835: data <= 'd3; 21836: data <= 'd6; 21837: data <= 'd6; 21838: data <= 'd6; 21839: data <= 'd6; 21840: data <= 'd6; 21841: data <= 'd6; 21842: data <= 'd6; 21843: data <= 'd3; 21844: data <= 'd2; 21845: data <= 'd0; 21846: data <= 'd0; 21847: data <= 'd0; 21848: data <= 'd0; 21849: data <= 'd0; 21850: data <= 'd0; 21851: data <= 'd0; 21852: data <= 'd0; 21853: data <= 'd0; 21854: data <= 'd0; 21855: data <= 'd0; 21856: data <= 'd0; 21857: data <= 'd0; 21858: data <= 'd0; 21859: data <= 'd0; 21860: data <= 'd0; 21861: data <= 'd0; 21862: data <= 'd0; 21863: data <= 'd0; 21864: data <= 'd0; 21865: data <= 'd2; 21866: data <= 'd1; 21867: data <= 'd3; 21868: data <= 'd6; 21869: data <= 'd6; 21870: data <= 'd6; 21871: data <= 'd6; 21872: data <= 'd6; 21873: data <= 'd6; 21874: data <= 'd6; 21875: data <= 'd3; 21876: data <= 'd1; 21877: data <= 'd2; 21878: data <= 'd0; 21879: data <= 'd0; 21880: data <= 'd0; 21881: data <= 'd0; 21882: data <= 'd0; 21883: data <= 'd0; 21884: data <= 'd0; 21885: data <= 'd0; 21886: data <= 'd0; 21887: data <= 'd0; 21888: data <= 'd0; 21889: data <= 'd0; 21890: data <= 'd0; 21891: data <= 'd0; 21892: data <= 'd0; 21893: data <= 'd0; 21894: data <= 'd0; 21895: data <= 'd0; 21896: data <= 'd0; 21897: data <= 'd2; 21898: data <= 'd1; 21899: data <= 'd3; 21900: data <= 'd3; 21901: data <= 'd6; 21902: data <= 'd6; 21903: data <= 'd6; 21904: data <= 'd6; 21905: data <= 'd6; 21906: data <= 'd3; 21907: data <= 'd3; 21908: data <= 'd1; 21909: data <= 'd2; 21910: data <= 'd0; 21911: data <= 'd0; 21912: data <= 'd0; 21913: data <= 'd0; 21914: data <= 'd0; 21915: data <= 'd0; 21916: data <= 'd0; 21917: data <= 'd0; 21918: data <= 'd0; 21919: data <= 'd0; 21920: data <= 'd0; 21921: data <= 'd0; 21922: data <= 'd0; 21923: data <= 'd0; 21924: data <= 'd0; 21925: data <= 'd0; 21926: data <= 'd0; 21927: data <= 'd0; 21928: data <= 'd2; 21929: data <= 'd1; 21930: data <= 'd1; 21931: data <= 'd1; 21932: data <= 'd3; 21933: data <= 'd3; 21934: data <= 'd3; 21935: data <= 'd3; 21936: data <= 'd3; 21937: data <= 'd3; 21938: data <= 'd3; 21939: data <= 'd1; 21940: data <= 'd1; 21941: data <= 'd1; 21942: data <= 'd2; 21943: data <= 'd0; 21944: data <= 'd0; 21945: data <= 'd0; 21946: data <= 'd0; 21947: data <= 'd0; 21948: data <= 'd0; 21949: data <= 'd0; 21950: data <= 'd0; 21951: data <= 'd0; 21952: data <= 'd0; 21953: data <= 'd0; 21954: data <= 'd0; 21955: data <= 'd0; 21956: data <= 'd0; 21957: data <= 'd0; 21958: data <= 'd0; 21959: data <= 'd0; 21960: data <= 'd5; 21961: data <= 'd5; 21962: data <= 'd1; 21963: data <= 'd3; 21964: data <= 'd3; 21965: data <= 'd3; 21966: data <= 'd3; 21967: data <= 'd3; 21968: data <= 'd3; 21969: data <= 'd3; 21970: data <= 'd3; 21971: data <= 'd3; 21972: data <= 'd1; 21973: data <= 'd5; 21974: data <= 'd5; 21975: data <= 'd0; 21976: data <= 'd0; 21977: data <= 'd0; 21978: data <= 'd0; 21979: data <= 'd0; 21980: data <= 'd0; 21981: data <= 'd0; 21982: data <= 'd0; 21983: data <= 'd0; 21984: data <= 'd0; 21985: data <= 'd0; 21986: data <= 'd0; 21987: data <= 'd0; 21988: data <= 'd0; 21989: data <= 'd0; 21990: data <= 'd0; 21991: data <= 'd2; 21992: data <= 'd3; 21993: data <= 'd3; 21994: data <= 'd1; 21995: data <= 'd3; 21996: data <= 'd3; 21997: data <= 'd3; 21998: data <= 'd3; 21999: data <= 'd6; 22000: data <= 'd3; 22001: data <= 'd3; 22002: data <= 'd3; 22003: data <= 'd3; 22004: data <= 'd1; 22005: data <= 'd3; 22006: data <= 'd3; 22007: data <= 'd2; 22008: data <= 'd0; 22009: data <= 'd0; 22010: data <= 'd0; 22011: data <= 'd0; 22012: data <= 'd0; 22013: data <= 'd0; 22014: data <= 'd0; 22015: data <= 'd0; 22016: data <= 'd0; 22017: data <= 'd0; 22018: data <= 'd0; 22019: data <= 'd0; 22020: data <= 'd0; 22021: data <= 'd0; 22022: data <= 'd0; 22023: data <= 'd2; 22024: data <= 'd3; 22025: data <= 'd3; 22026: data <= 'd3; 22027: data <= 'd1; 22028: data <= 'd3; 22029: data <= 'd3; 22030: data <= 'd6; 22031: data <= 'd6; 22032: data <= 'd6; 22033: data <= 'd3; 22034: data <= 'd3; 22035: data <= 'd1; 22036: data <= 'd3; 22037: data <= 'd3; 22038: data <= 'd3; 22039: data <= 'd2; 22040: data <= 'd0; 22041: data <= 'd0; 22042: data <= 'd0; 22043: data <= 'd0; 22044: data <= 'd0; 22045: data <= 'd0; 22046: data <= 'd0; 22047: data <= 'd0; 22048: data <= 'd0; 22049: data <= 'd0; 22050: data <= 'd0; 22051: data <= 'd0; 22052: data <= 'd0; 22053: data <= 'd0; 22054: data <= 'd0; 22055: data <= 'd2; 22056: data <= 'd1; 22057: data <= 'd1; 22058: data <= 'd3; 22059: data <= 'd1; 22060: data <= 'd5; 22061: data <= 'd3; 22062: data <= 'd6; 22063: data <= 'd6; 22064: data <= 'd6; 22065: data <= 'd3; 22066: data <= 'd5; 22067: data <= 'd1; 22068: data <= 'd3; 22069: data <= 'd1; 22070: data <= 'd1; 22071: data <= 'd2; 22072: data <= 'd0; 22073: data <= 'd0; 22074: data <= 'd0; 22075: data <= 'd0; 22076: data <= 'd0; 22077: data <= 'd0; 22078: data <= 'd0; 22079: data <= 'd0; 22080: data <= 'd0; 22081: data <= 'd0; 22082: data <= 'd0; 22083: data <= 'd0; 22084: data <= 'd0; 22085: data <= 'd0; 22086: data <= 'd0; 22087: data <= 'd0; 22088: data <= 'd2; 22089: data <= 'd2; 22090: data <= 'd1; 22091: data <= 'd1; 22092: data <= 'd5; 22093: data <= 'd3; 22094: data <= 'd3; 22095: data <= 'd6; 22096: data <= 'd3; 22097: data <= 'd3; 22098: data <= 'd5; 22099: data <= 'd1; 22100: data <= 'd1; 22101: data <= 'd2; 22102: data <= 'd2; 22103: data <= 'd0; 22104: data <= 'd0; 22105: data <= 'd0; 22106: data <= 'd0; 22107: data <= 'd0; 22108: data <= 'd0; 22109: data <= 'd0; 22110: data <= 'd0; 22111: data <= 'd0; 22112: data <= 'd0; 22113: data <= 'd0; 22114: data <= 'd0; 22115: data <= 'd0; 22116: data <= 'd0; 22117: data <= 'd0; 22118: data <= 'd0; 22119: data <= 'd0; 22120: data <= 'd2; 22121: data <= 'd8; 22122: data <= 'd2; 22123: data <= 'd2; 22124: data <= 'd2; 22125: data <= 'd1; 22126: data <= 'd3; 22127: data <= 'd3; 22128: data <= 'd3; 22129: data <= 'd1; 22130: data <= 'd2; 22131: data <= 'd2; 22132: data <= 'd2; 22133: data <= 'd8; 22134: data <= 'd2; 22135: data <= 'd0; 22136: data <= 'd0; 22137: data <= 'd0; 22138: data <= 'd0; 22139: data <= 'd0; 22140: data <= 'd0; 22141: data <= 'd0; 22142: data <= 'd0; 22143: data <= 'd0; 22144: data <= 'd0; 22145: data <= 'd0; 22146: data <= 'd0; 22147: data <= 'd0; 22148: data <= 'd0; 22149: data <= 'd0; 22150: data <= 'd0; 22151: data <= 'd0; 22152: data <= 'd0; 22153: data <= 'd2; 22154: data <= 'd8; 22155: data <= 'd8; 22156: data <= 'd8; 22157: data <= 'd2; 22158: data <= 'd3; 22159: data <= 'd3; 22160: data <= 'd3; 22161: data <= 'd1; 22162: data <= 'd2; 22163: data <= 'd8; 22164: data <= 'd8; 22165: data <= 'd2; 22166: data <= 'd0; 22167: data <= 'd0; 22168: data <= 'd0; 22169: data <= 'd0; 22170: data <= 'd0; 22171: data <= 'd0; 22172: data <= 'd0; 22173: data <= 'd0; 22174: data <= 'd0; 22175: data <= 'd0; 22176: data <= 'd0; 22177: data <= 'd0; 22178: data <= 'd0; 22179: data <= 'd0; 22180: data <= 'd0; 22181: data <= 'd0; 22182: data <= 'd0; 22183: data <= 'd0; 22184: data <= 'd2; 22185: data <= 'd9; 22186: data <= 'd5; 22187: data <= 'd8; 22188: data <= 'd9; 22189: data <= 'd8; 22190: data <= 'd2; 22191: data <= 'd1; 22192: data <= 'd3; 22193: data <= 'd1; 22194: data <= 'd2; 22195: data <= 'd8; 22196: data <= 'd9; 22197: data <= 'd2; 22198: data <= 'd0; 22199: data <= 'd0; 22200: data <= 'd0; 22201: data <= 'd0; 22202: data <= 'd0; 22203: data <= 'd0; 22204: data <= 'd0; 22205: data <= 'd0; 22206: data <= 'd0; 22207: data <= 'd0; 22208: data <= 'd0; 22209: data <= 'd0; 22210: data <= 'd0; 22211: data <= 'd0; 22212: data <= 'd0; 22213: data <= 'd0; 22214: data <= 'd0; 22215: data <= 'd0; 22216: data <= 'd2; 22217: data <= 'd9; 22218: data <= 'd4; 22219: data <= 'd9; 22220: data <= 'd9; 22221: data <= 'd9; 22222: data <= 'd8; 22223: data <= 'd2; 22224: data <= 'd2; 22225: data <= 'd2; 22226: data <= 'd8; 22227: data <= 'd8; 22228: data <= 'd2; 22229: data <= 'd2; 22230: data <= 'd0; 22231: data <= 'd0; 22232: data <= 'd0; 22233: data <= 'd0; 22234: data <= 'd0; 22235: data <= 'd0; 22236: data <= 'd0; 22237: data <= 'd0; 22238: data <= 'd0; 22239: data <= 'd0; 22240: data <= 'd0; 22241: data <= 'd0; 22242: data <= 'd0; 22243: data <= 'd0; 22244: data <= 'd0; 22245: data <= 'd0; 22246: data <= 'd0; 22247: data <= 'd0; 22248: data <= 'd0; 22249: data <= 'd2; 22250: data <= 'd7; 22251: data <= 'd1; 22252: data <= 'd3; 22253: data <= 'd3; 22254: data <= 'd3; 22255: data <= 'd1; 22256: data <= 'd1; 22257: data <= 'd1; 22258: data <= 'd3; 22259: data <= 'd1; 22260: data <= 'd7; 22261: data <= 'd2; 22262: data <= 'd0; 22263: data <= 'd0; 22264: data <= 'd0; 22265: data <= 'd0; 22266: data <= 'd0; 22267: data <= 'd0; 22268: data <= 'd0; 22269: data <= 'd0; 22270: data <= 'd0; 22271: data <= 'd0; 22272: data <= 'd0; 22273: data <= 'd0; 22274: data <= 'd0; 22275: data <= 'd0; 22276: data <= 'd0; 22277: data <= 'd0; 22278: data <= 'd0; 22279: data <= 'd0; 22280: data <= 'd0; 22281: data <= 'd2; 22282: data <= 'd7; 22283: data <= 'd5; 22284: data <= 'd3; 22285: data <= 'd3; 22286: data <= 'd3; 22287: data <= 'd3; 22288: data <= 'd3; 22289: data <= 'd3; 22290: data <= 'd3; 22291: data <= 'd5; 22292: data <= 'd7; 22293: data <= 'd4; 22294: data <= 'd2; 22295: data <= 'd0; 22296: data <= 'd0; 22297: data <= 'd0; 22298: data <= 'd0; 22299: data <= 'd0; 22300: data <= 'd0; 22301: data <= 'd0; 22302: data <= 'd0; 22303: data <= 'd0; 22304: data <= 'd0; 22305: data <= 'd0; 22306: data <= 'd0; 22307: data <= 'd0; 22308: data <= 'd0; 22309: data <= 'd0; 22310: data <= 'd0; 22311: data <= 'd0; 22312: data <= 'd0; 22313: data <= 'd0; 22314: data <= 'd2; 22315: data <= 'd1; 22316: data <= 'd3; 22317: data <= 'd3; 22318: data <= 'd3; 22319: data <= 'd3; 22320: data <= 'd3; 22321: data <= 'd3; 22322: data <= 'd3; 22323: data <= 'd1; 22324: data <= 'd4; 22325: data <= 'd9; 22326: data <= 'd2; 22327: data <= 'd0; 22328: data <= 'd0; 22329: data <= 'd0; 22330: data <= 'd0; 22331: data <= 'd0; 22332: data <= 'd0; 22333: data <= 'd0; 22334: data <= 'd0; 22335: data <= 'd0; 22336: data <= 'd0; 22337: data <= 'd0; 22338: data <= 'd0; 22339: data <= 'd0; 22340: data <= 'd0; 22341: data <= 'd0; 22342: data <= 'd0; 22343: data <= 'd0; 22344: data <= 'd0; 22345: data <= 'd0; 22346: data <= 'd2; 22347: data <= 'd1; 22348: data <= 'd1; 22349: data <= 'd3; 22350: data <= 'd3; 22351: data <= 'd3; 22352: data <= 'd3; 22353: data <= 'd3; 22354: data <= 'd1; 22355: data <= 'd1; 22356: data <= 'd2; 22357: data <= 'd9; 22358: data <= 'd2; 22359: data <= 'd0; 22360: data <= 'd0; 22361: data <= 'd0; 22362: data <= 'd0; 22363: data <= 'd0; 22364: data <= 'd0; 22365: data <= 'd0; 22366: data <= 'd0; 22367: data <= 'd0; 22368: data <= 'd0; 22369: data <= 'd0; 22370: data <= 'd0; 22371: data <= 'd0; 22372: data <= 'd0; 22373: data <= 'd0; 22374: data <= 'd0; 22375: data <= 'd0; 22376: data <= 'd0; 22377: data <= 'd0; 22378: data <= 'd2; 22379: data <= 'd2; 22380: data <= 'd2; 22381: data <= 'd2; 22382: data <= 'd5; 22383: data <= 'd5; 22384: data <= 'd5; 22385: data <= 'd2; 22386: data <= 'd2; 22387: data <= 'd2; 22388: data <= 'd2; 22389: data <= 'd2; 22390: data <= 'd0; 22391: data <= 'd0; 22392: data <= 'd0; 22393: data <= 'd0; 22394: data <= 'd0; 22395: data <= 'd0; 22396: data <= 'd0; 22397: data <= 'd0; 22398: data <= 'd0; 22399: data <= 'd0; 22400: data <= 'd0; 22401: data <= 'd0; 22402: data <= 'd0; 22403: data <= 'd0; 22404: data <= 'd0; 22405: data <= 'd0; 22406: data <= 'd0; 22407: data <= 'd0; 22408: data <= 'd0; 22409: data <= 'd0; 22410: data <= 'd2; 22411: data <= 'd1; 22412: data <= 'd1; 22413: data <= 'd3; 22414: data <= 'd3; 22415: data <= 'd3; 22416: data <= 'd3; 22417: data <= 'd3; 22418: data <= 'd1; 22419: data <= 'd1; 22420: data <= 'd2; 22421: data <= 'd0; 22422: data <= 'd0; 22423: data <= 'd0; 22424: data <= 'd0; 22425: data <= 'd0; 22426: data <= 'd0; 22427: data <= 'd0; 22428: data <= 'd0; 22429: data <= 'd0; 22430: data <= 'd0; 22431: data <= 'd0; 22432: data <= 'd0; 22433: data <= 'd0; 22434: data <= 'd0; 22435: data <= 'd0; 22436: data <= 'd0; 22437: data <= 'd0; 22438: data <= 'd0; 22439: data <= 'd0; 22440: data <= 'd0; 22441: data <= 'd0; 22442: data <= 'd2; 22443: data <= 'd7; 22444: data <= 'd7; 22445: data <= 'd4; 22446: data <= 'd2; 22447: data <= 'd2; 22448: data <= 'd2; 22449: data <= 'd2; 22450: data <= 'd7; 22451: data <= 'd7; 22452: data <= 'd2; 22453: data <= 'd0; 22454: data <= 'd0; 22455: data <= 'd0; 22456: data <= 'd0; 22457: data <= 'd0; 22458: data <= 'd0; 22459: data <= 'd0; 22460: data <= 'd0; 22461: data <= 'd0; 22462: data <= 'd0; 22463: data <= 'd0; 22464: data <= 'd0; 22465: data <= 'd0; 22466: data <= 'd0; 22467: data <= 'd0; 22468: data <= 'd0; 22469: data <= 'd0; 22470: data <= 'd0; 22471: data <= 'd0; 22472: data <= 'd0; 22473: data <= 'd0; 22474: data <= 'd2; 22475: data <= 'd4; 22476: data <= 'd7; 22477: data <= 'd2; 22478: data <= 'd0; 22479: data <= 'd0; 22480: data <= 'd0; 22481: data <= 'd0; 22482: data <= 'd2; 22483: data <= 'd2; 22484: data <= 'd2; 22485: data <= 'd0; 22486: data <= 'd0; 22487: data <= 'd0; 22488: data <= 'd0; 22489: data <= 'd0; 22490: data <= 'd0; 22491: data <= 'd0; 22492: data <= 'd0; 22493: data <= 'd0; 22494: data <= 'd0; 22495: data <= 'd0; 22496: data <= 'd0; 22497: data <= 'd0; 22498: data <= 'd0; 22499: data <= 'd0; 22500: data <= 'd0; 22501: data <= 'd0; 22502: data <= 'd0; 22503: data <= 'd0; 22504: data <= 'd0; 22505: data <= 'd0; 22506: data <= 'd0; 22507: data <= 'd2; 22508: data <= 'd2; 22509: data <= 'd2; 22510: data <= 'd0; 22511: data <= 'd0; 22512: data <= 'd0; 22513: data <= 'd0; 22514: data <= 'd0; 22515: data <= 'd0; 22516: data <= 'd0; 22517: data <= 'd0; 22518: data <= 'd0; 22519: data <= 'd0; 22520: data <= 'd0; 22521: data <= 'd0; 22522: data <= 'd0; 22523: data <= 'd0; 22524: data <= 'd0; 22525: data <= 'd0; 22526: data <= 'd0; 22527: data <= 'd0; 22528: data <= 'd0; 22529: data <= 'd0; 22530: data <= 'd0; 22531: data <= 'd0; 22532: data <= 'd0; 22533: data <= 'd0; 22534: data <= 'd0; 22535: data <= 'd0; 22536: data <= 'd0; 22537: data <= 'd0; 22538: data <= 'd0; 22539: data <= 'd0; 22540: data <= 'd0; 22541: data <= 'd0; 22542: data <= 'd0; 22543: data <= 'd0; 22544: data <= 'd0; 22545: data <= 'd0; 22546: data <= 'd0; 22547: data <= 'd0; 22548: data <= 'd0; 22549: data <= 'd0; 22550: data <= 'd0; 22551: data <= 'd0; 22552: data <= 'd0; 22553: data <= 'd0; 22554: data <= 'd0; 22555: data <= 'd0; 22556: data <= 'd0; 22557: data <= 'd0; 22558: data <= 'd0; 22559: data <= 'd0; 22560: data <= 'd0; 22561: data <= 'd0; 22562: data <= 'd0; 22563: data <= 'd0; 22564: data <= 'd0; 22565: data <= 'd0; 22566: data <= 'd0; 22567: data <= 'd0; 22568: data <= 'd0; 22569: data <= 'd0; 22570: data <= 'd0; 22571: data <= 'd0; 22572: data <= 'd0; 22573: data <= 'd0; 22574: data <= 'd0; 22575: data <= 'd0; 22576: data <= 'd0; 22577: data <= 'd0; 22578: data <= 'd0; 22579: data <= 'd0; 22580: data <= 'd0; 22581: data <= 'd0; 22582: data <= 'd0; 22583: data <= 'd0; 22584: data <= 'd0; 22585: data <= 'd0; 22586: data <= 'd0; 22587: data <= 'd0; 22588: data <= 'd0; 22589: data <= 'd0; 22590: data <= 'd0; 22591: data <= 'd0; 22592: data <= 'd0; 22593: data <= 'd0; 22594: data <= 'd0; 22595: data <= 'd0; 22596: data <= 'd0; 22597: data <= 'd0; 22598: data <= 'd0; 22599: data <= 'd0; 22600: data <= 'd0; 22601: data <= 'd0; 22602: data <= 'd0; 22603: data <= 'd0; 22604: data <= 'd0; 22605: data <= 'd0; 22606: data <= 'd0; 22607: data <= 'd0; 22608: data <= 'd0; 22609: data <= 'd0; 22610: data <= 'd0; 22611: data <= 'd0; 22612: data <= 'd0; 22613: data <= 'd0; 22614: data <= 'd0; 22615: data <= 'd0; 22616: data <= 'd0; 22617: data <= 'd0; 22618: data <= 'd0; 22619: data <= 'd0; 22620: data <= 'd0; 22621: data <= 'd0; 22622: data <= 'd0; 22623: data <= 'd0; 22624: data <= 'd0; 22625: data <= 'd0; 22626: data <= 'd0; 22627: data <= 'd0; 22628: data <= 'd0; 22629: data <= 'd0; 22630: data <= 'd0; 22631: data <= 'd0; 22632: data <= 'd0; 22633: data <= 'd0; 22634: data <= 'd0; 22635: data <= 'd0; 22636: data <= 'd0; 22637: data <= 'd0; 22638: data <= 'd0; 22639: data <= 'd0; 22640: data <= 'd0; 22641: data <= 'd0; 22642: data <= 'd0; 22643: data <= 'd0; 22644: data <= 'd0; 22645: data <= 'd0; 22646: data <= 'd0; 22647: data <= 'd0; 22648: data <= 'd0; 22649: data <= 'd0; 22650: data <= 'd0; 22651: data <= 'd0; 22652: data <= 'd0; 22653: data <= 'd0; 22654: data <= 'd0; 22655: data <= 'd0; 22656: data <= 'd0; 22657: data <= 'd0; 22658: data <= 'd0; 22659: data <= 'd0; 22660: data <= 'd0; 22661: data <= 'd0; 22662: data <= 'd0; 22663: data <= 'd0; 22664: data <= 'd0; 22665: data <= 'd0; 22666: data <= 'd0; 22667: data <= 'd0; 22668: data <= 'd0; 22669: data <= 'd0; 22670: data <= 'd0; 22671: data <= 'd0; 22672: data <= 'd0; 22673: data <= 'd0; 22674: data <= 'd0; 22675: data <= 'd0; 22676: data <= 'd0; 22677: data <= 'd0; 22678: data <= 'd0; 22679: data <= 'd0; 22680: data <= 'd0; 22681: data <= 'd0; 22682: data <= 'd0; 22683: data <= 'd0; 22684: data <= 'd0; 22685: data <= 'd0; 22686: data <= 'd0; 22687: data <= 'd0; 22688: data <= 'd0; 22689: data <= 'd0; 22690: data <= 'd0; 22691: data <= 'd0; 22692: data <= 'd0; 22693: data <= 'd0; 22694: data <= 'd0; 22695: data <= 'd0; 22696: data <= 'd0; 22697: data <= 'd0; 22698: data <= 'd0; 22699: data <= 'd0; 22700: data <= 'd0; 22701: data <= 'd0; 22702: data <= 'd0; 22703: data <= 'd0; 22704: data <= 'd0; 22705: data <= 'd0; 22706: data <= 'd0; 22707: data <= 'd0; 22708: data <= 'd0; 22709: data <= 'd0; 22710: data <= 'd0; 22711: data <= 'd0; 22712: data <= 'd0; 22713: data <= 'd0; 22714: data <= 'd0; 22715: data <= 'd0; 22716: data <= 'd0; 22717: data <= 'd0; 22718: data <= 'd0; 22719: data <= 'd0; 22720: data <= 'd0; 22721: data <= 'd0; 22722: data <= 'd0; 22723: data <= 'd0; 22724: data <= 'd0; 22725: data <= 'd0; 22726: data <= 'd0; 22727: data <= 'd0; 22728: data <= 'd0; 22729: data <= 'd0; 22730: data <= 'd0; 22731: data <= 'd0; 22732: data <= 'd0; 22733: data <= 'd0; 22734: data <= 'd0; 22735: data <= 'd0; 22736: data <= 'd0; 22737: data <= 'd0; 22738: data <= 'd0; 22739: data <= 'd0; 22740: data <= 'd0; 22741: data <= 'd0; 22742: data <= 'd0; 22743: data <= 'd0; 22744: data <= 'd0; 22745: data <= 'd0; 22746: data <= 'd0; 22747: data <= 'd0; 22748: data <= 'd0; 22749: data <= 'd0; 22750: data <= 'd0; 22751: data <= 'd0; 22752: data <= 'd0; 22753: data <= 'd0; 22754: data <= 'd0; 22755: data <= 'd0; 22756: data <= 'd0; 22757: data <= 'd0; 22758: data <= 'd0; 22759: data <= 'd0; 22760: data <= 'd0; 22761: data <= 'd0; 22762: data <= 'd0; 22763: data <= 'd0; 22764: data <= 'd0; 22765: data <= 'd0; 22766: data <= 'd0; 22767: data <= 'd0; 22768: data <= 'd0; 22769: data <= 'd0; 22770: data <= 'd0; 22771: data <= 'd0; 22772: data <= 'd0; 22773: data <= 'd0; 22774: data <= 'd0; 22775: data <= 'd0; 22776: data <= 'd0; 22777: data <= 'd0; 22778: data <= 'd0; 22779: data <= 'd0; 22780: data <= 'd0; 22781: data <= 'd0; 22782: data <= 'd0; 22783: data <= 'd0; 22784: data <= 'd0; 22785: data <= 'd0; 22786: data <= 'd0; 22787: data <= 'd0; 22788: data <= 'd0; 22789: data <= 'd0; 22790: data <= 'd0; 22791: data <= 'd0; 22792: data <= 'd0; 22793: data <= 'd0; 22794: data <= 'd0; 22795: data <= 'd0; 22796: data <= 'd0; 22797: data <= 'd2; 22798: data <= 'd2; 22799: data <= 'd2; 22800: data <= 'd2; 22801: data <= 'd2; 22802: data <= 'd0; 22803: data <= 'd0; 22804: data <= 'd0; 22805: data <= 'd0; 22806: data <= 'd0; 22807: data <= 'd0; 22808: data <= 'd0; 22809: data <= 'd0; 22810: data <= 'd0; 22811: data <= 'd0; 22812: data <= 'd0; 22813: data <= 'd0; 22814: data <= 'd0; 22815: data <= 'd0; 22816: data <= 'd0; 22817: data <= 'd0; 22818: data <= 'd0; 22819: data <= 'd0; 22820: data <= 'd0; 22821: data <= 'd0; 22822: data <= 'd0; 22823: data <= 'd0; 22824: data <= 'd0; 22825: data <= 'd0; 22826: data <= 'd0; 22827: data <= 'd2; 22828: data <= 'd2; 22829: data <= 'd6; 22830: data <= 'd6; 22831: data <= 'd6; 22832: data <= 'd6; 22833: data <= 'd6; 22834: data <= 'd2; 22835: data <= 'd2; 22836: data <= 'd0; 22837: data <= 'd0; 22838: data <= 'd0; 22839: data <= 'd0; 22840: data <= 'd0; 22841: data <= 'd0; 22842: data <= 'd0; 22843: data <= 'd0; 22844: data <= 'd0; 22845: data <= 'd0; 22846: data <= 'd0; 22847: data <= 'd0; 22848: data <= 'd0; 22849: data <= 'd0; 22850: data <= 'd0; 22851: data <= 'd0; 22852: data <= 'd0; 22853: data <= 'd0; 22854: data <= 'd0; 22855: data <= 'd0; 22856: data <= 'd0; 22857: data <= 'd0; 22858: data <= 'd2; 22859: data <= 'd3; 22860: data <= 'd6; 22861: data <= 'd6; 22862: data <= 'd6; 22863: data <= 'd6; 22864: data <= 'd6; 22865: data <= 'd6; 22866: data <= 'd6; 22867: data <= 'd3; 22868: data <= 'd2; 22869: data <= 'd0; 22870: data <= 'd0; 22871: data <= 'd0; 22872: data <= 'd0; 22873: data <= 'd0; 22874: data <= 'd0; 22875: data <= 'd0; 22876: data <= 'd0; 22877: data <= 'd0; 22878: data <= 'd0; 22879: data <= 'd0; 22880: data <= 'd0; 22881: data <= 'd0; 22882: data <= 'd0; 22883: data <= 'd0; 22884: data <= 'd0; 22885: data <= 'd0; 22886: data <= 'd0; 22887: data <= 'd0; 22888: data <= 'd0; 22889: data <= 'd2; 22890: data <= 'd1; 22891: data <= 'd3; 22892: data <= 'd6; 22893: data <= 'd6; 22894: data <= 'd6; 22895: data <= 'd6; 22896: data <= 'd6; 22897: data <= 'd6; 22898: data <= 'd6; 22899: data <= 'd3; 22900: data <= 'd1; 22901: data <= 'd2; 22902: data <= 'd0; 22903: data <= 'd0; 22904: data <= 'd0; 22905: data <= 'd0; 22906: data <= 'd0; 22907: data <= 'd0; 22908: data <= 'd0; 22909: data <= 'd0; 22910: data <= 'd0; 22911: data <= 'd0; 22912: data <= 'd0; 22913: data <= 'd0; 22914: data <= 'd0; 22915: data <= 'd0; 22916: data <= 'd0; 22917: data <= 'd0; 22918: data <= 'd0; 22919: data <= 'd0; 22920: data <= 'd0; 22921: data <= 'd2; 22922: data <= 'd1; 22923: data <= 'd3; 22924: data <= 'd3; 22925: data <= 'd6; 22926: data <= 'd6; 22927: data <= 'd6; 22928: data <= 'd6; 22929: data <= 'd6; 22930: data <= 'd3; 22931: data <= 'd3; 22932: data <= 'd1; 22933: data <= 'd2; 22934: data <= 'd0; 22935: data <= 'd0; 22936: data <= 'd0; 22937: data <= 'd0; 22938: data <= 'd0; 22939: data <= 'd0; 22940: data <= 'd0; 22941: data <= 'd0; 22942: data <= 'd0; 22943: data <= 'd0; 22944: data <= 'd0; 22945: data <= 'd0; 22946: data <= 'd0; 22947: data <= 'd0; 22948: data <= 'd0; 22949: data <= 'd0; 22950: data <= 'd0; 22951: data <= 'd0; 22952: data <= 'd2; 22953: data <= 'd1; 22954: data <= 'd1; 22955: data <= 'd1; 22956: data <= 'd3; 22957: data <= 'd3; 22958: data <= 'd3; 22959: data <= 'd3; 22960: data <= 'd3; 22961: data <= 'd3; 22962: data <= 'd3; 22963: data <= 'd1; 22964: data <= 'd1; 22965: data <= 'd1; 22966: data <= 'd2; 22967: data <= 'd0; 22968: data <= 'd0; 22969: data <= 'd0; 22970: data <= 'd0; 22971: data <= 'd0; 22972: data <= 'd0; 22973: data <= 'd0; 22974: data <= 'd0; 22975: data <= 'd0; 22976: data <= 'd0; 22977: data <= 'd0; 22978: data <= 'd0; 22979: data <= 'd0; 22980: data <= 'd0; 22981: data <= 'd0; 22982: data <= 'd0; 22983: data <= 'd0; 22984: data <= 'd5; 22985: data <= 'd5; 22986: data <= 'd1; 22987: data <= 'd3; 22988: data <= 'd3; 22989: data <= 'd3; 22990: data <= 'd3; 22991: data <= 'd3; 22992: data <= 'd3; 22993: data <= 'd3; 22994: data <= 'd3; 22995: data <= 'd3; 22996: data <= 'd1; 22997: data <= 'd5; 22998: data <= 'd5; 22999: data <= 'd0; 23000: data <= 'd0; 23001: data <= 'd0; 23002: data <= 'd0; 23003: data <= 'd0; 23004: data <= 'd0; 23005: data <= 'd0; 23006: data <= 'd0; 23007: data <= 'd0; 23008: data <= 'd0; 23009: data <= 'd0; 23010: data <= 'd0; 23011: data <= 'd0; 23012: data <= 'd0; 23013: data <= 'd0; 23014: data <= 'd0; 23015: data <= 'd2; 23016: data <= 'd3; 23017: data <= 'd3; 23018: data <= 'd1; 23019: data <= 'd3; 23020: data <= 'd3; 23021: data <= 'd3; 23022: data <= 'd3; 23023: data <= 'd6; 23024: data <= 'd3; 23025: data <= 'd3; 23026: data <= 'd3; 23027: data <= 'd3; 23028: data <= 'd1; 23029: data <= 'd3; 23030: data <= 'd3; 23031: data <= 'd2; 23032: data <= 'd0; 23033: data <= 'd0; 23034: data <= 'd0; 23035: data <= 'd0; 23036: data <= 'd0; 23037: data <= 'd0; 23038: data <= 'd0; 23039: data <= 'd0; 23040: data <= 'd0; 23041: data <= 'd0; 23042: data <= 'd0; 23043: data <= 'd0; 23044: data <= 'd0; 23045: data <= 'd0; 23046: data <= 'd0; 23047: data <= 'd2; 23048: data <= 'd3; 23049: data <= 'd3; 23050: data <= 'd3; 23051: data <= 'd1; 23052: data <= 'd3; 23053: data <= 'd3; 23054: data <= 'd6; 23055: data <= 'd6; 23056: data <= 'd6; 23057: data <= 'd3; 23058: data <= 'd3; 23059: data <= 'd1; 23060: data <= 'd3; 23061: data <= 'd3; 23062: data <= 'd3; 23063: data <= 'd2; 23064: data <= 'd0; 23065: data <= 'd0; 23066: data <= 'd0; 23067: data <= 'd0; 23068: data <= 'd0; 23069: data <= 'd0; 23070: data <= 'd0; 23071: data <= 'd0; 23072: data <= 'd0; 23073: data <= 'd0; 23074: data <= 'd0; 23075: data <= 'd0; 23076: data <= 'd0; 23077: data <= 'd0; 23078: data <= 'd0; 23079: data <= 'd2; 23080: data <= 'd1; 23081: data <= 'd1; 23082: data <= 'd3; 23083: data <= 'd1; 23084: data <= 'd5; 23085: data <= 'd3; 23086: data <= 'd6; 23087: data <= 'd6; 23088: data <= 'd6; 23089: data <= 'd3; 23090: data <= 'd5; 23091: data <= 'd1; 23092: data <= 'd3; 23093: data <= 'd1; 23094: data <= 'd1; 23095: data <= 'd2; 23096: data <= 'd0; 23097: data <= 'd0; 23098: data <= 'd0; 23099: data <= 'd0; 23100: data <= 'd0; 23101: data <= 'd0; 23102: data <= 'd0; 23103: data <= 'd0; 23104: data <= 'd0; 23105: data <= 'd0; 23106: data <= 'd0; 23107: data <= 'd0; 23108: data <= 'd0; 23109: data <= 'd0; 23110: data <= 'd0; 23111: data <= 'd0; 23112: data <= 'd2; 23113: data <= 'd2; 23114: data <= 'd1; 23115: data <= 'd1; 23116: data <= 'd5; 23117: data <= 'd3; 23118: data <= 'd3; 23119: data <= 'd6; 23120: data <= 'd3; 23121: data <= 'd3; 23122: data <= 'd5; 23123: data <= 'd1; 23124: data <= 'd1; 23125: data <= 'd2; 23126: data <= 'd2; 23127: data <= 'd0; 23128: data <= 'd0; 23129: data <= 'd0; 23130: data <= 'd0; 23131: data <= 'd0; 23132: data <= 'd0; 23133: data <= 'd0; 23134: data <= 'd0; 23135: data <= 'd0; 23136: data <= 'd0; 23137: data <= 'd0; 23138: data <= 'd0; 23139: data <= 'd0; 23140: data <= 'd0; 23141: data <= 'd0; 23142: data <= 'd0; 23143: data <= 'd0; 23144: data <= 'd2; 23145: data <= 'd8; 23146: data <= 'd2; 23147: data <= 'd2; 23148: data <= 'd2; 23149: data <= 'd1; 23150: data <= 'd3; 23151: data <= 'd3; 23152: data <= 'd3; 23153: data <= 'd1; 23154: data <= 'd2; 23155: data <= 'd2; 23156: data <= 'd2; 23157: data <= 'd8; 23158: data <= 'd2; 23159: data <= 'd0; 23160: data <= 'd0; 23161: data <= 'd0; 23162: data <= 'd0; 23163: data <= 'd0; 23164: data <= 'd0; 23165: data <= 'd0; 23166: data <= 'd0; 23167: data <= 'd0; 23168: data <= 'd0; 23169: data <= 'd0; 23170: data <= 'd0; 23171: data <= 'd0; 23172: data <= 'd0; 23173: data <= 'd0; 23174: data <= 'd0; 23175: data <= 'd0; 23176: data <= 'd0; 23177: data <= 'd2; 23178: data <= 'd8; 23179: data <= 'd8; 23180: data <= 'd2; 23181: data <= 'd1; 23182: data <= 'd3; 23183: data <= 'd3; 23184: data <= 'd3; 23185: data <= 'd1; 23186: data <= 'd2; 23187: data <= 'd8; 23188: data <= 'd8; 23189: data <= 'd2; 23190: data <= 'd0; 23191: data <= 'd0; 23192: data <= 'd0; 23193: data <= 'd0; 23194: data <= 'd0; 23195: data <= 'd0; 23196: data <= 'd0; 23197: data <= 'd0; 23198: data <= 'd0; 23199: data <= 'd0; 23200: data <= 'd0; 23201: data <= 'd0; 23202: data <= 'd0; 23203: data <= 'd0; 23204: data <= 'd0; 23205: data <= 'd0; 23206: data <= 'd0; 23207: data <= 'd0; 23208: data <= 'd0; 23209: data <= 'd2; 23210: data <= 'd9; 23211: data <= 'd8; 23212: data <= 'd8; 23213: data <= 'd2; 23214: data <= 'd1; 23215: data <= 'd3; 23216: data <= 'd1; 23217: data <= 'd2; 23218: data <= 'd8; 23219: data <= 'd8; 23220: data <= 'd9; 23221: data <= 'd2; 23222: data <= 'd0; 23223: data <= 'd0; 23224: data <= 'd0; 23225: data <= 'd0; 23226: data <= 'd0; 23227: data <= 'd0; 23228: data <= 'd0; 23229: data <= 'd0; 23230: data <= 'd0; 23231: data <= 'd0; 23232: data <= 'd0; 23233: data <= 'd0; 23234: data <= 'd0; 23235: data <= 'd0; 23236: data <= 'd0; 23237: data <= 'd0; 23238: data <= 'd0; 23239: data <= 'd0; 23240: data <= 'd0; 23241: data <= 'd2; 23242: data <= 'd2; 23243: data <= 'd8; 23244: data <= 'd8; 23245: data <= 'd8; 23246: data <= 'd2; 23247: data <= 'd2; 23248: data <= 'd2; 23249: data <= 'd8; 23250: data <= 'd8; 23251: data <= 'd9; 23252: data <= 'd8; 23253: data <= 'd2; 23254: data <= 'd0; 23255: data <= 'd0; 23256: data <= 'd0; 23257: data <= 'd0; 23258: data <= 'd0; 23259: data <= 'd0; 23260: data <= 'd0; 23261: data <= 'd0; 23262: data <= 'd0; 23263: data <= 'd0; 23264: data <= 'd0; 23265: data <= 'd0; 23266: data <= 'd0; 23267: data <= 'd0; 23268: data <= 'd0; 23269: data <= 'd0; 23270: data <= 'd0; 23271: data <= 'd0; 23272: data <= 'd0; 23273: data <= 'd2; 23274: data <= 'd7; 23275: data <= 'd1; 23276: data <= 'd3; 23277: data <= 'd3; 23278: data <= 'd1; 23279: data <= 'd1; 23280: data <= 'd1; 23281: data <= 'd3; 23282: data <= 'd3; 23283: data <= 'd1; 23284: data <= 'd7; 23285: data <= 'd2; 23286: data <= 'd0; 23287: data <= 'd0; 23288: data <= 'd0; 23289: data <= 'd0; 23290: data <= 'd0; 23291: data <= 'd0; 23292: data <= 'd0; 23293: data <= 'd0; 23294: data <= 'd0; 23295: data <= 'd0; 23296: data <= 'd0; 23297: data <= 'd0; 23298: data <= 'd0; 23299: data <= 'd0; 23300: data <= 'd0; 23301: data <= 'd0; 23302: data <= 'd0; 23303: data <= 'd0; 23304: data <= 'd2; 23305: data <= 'd7; 23306: data <= 'd7; 23307: data <= 'd5; 23308: data <= 'd3; 23309: data <= 'd3; 23310: data <= 'd3; 23311: data <= 'd3; 23312: data <= 'd3; 23313: data <= 'd3; 23314: data <= 'd3; 23315: data <= 'd5; 23316: data <= 'd7; 23317: data <= 'd7; 23318: data <= 'd2; 23319: data <= 'd0; 23320: data <= 'd0; 23321: data <= 'd0; 23322: data <= 'd0; 23323: data <= 'd0; 23324: data <= 'd0; 23325: data <= 'd0; 23326: data <= 'd0; 23327: data <= 'd0; 23328: data <= 'd0; 23329: data <= 'd0; 23330: data <= 'd0; 23331: data <= 'd0; 23332: data <= 'd0; 23333: data <= 'd0; 23334: data <= 'd0; 23335: data <= 'd0; 23336: data <= 'd2; 23337: data <= 'd4; 23338: data <= 'd1; 23339: data <= 'd1; 23340: data <= 'd3; 23341: data <= 'd3; 23342: data <= 'd3; 23343: data <= 'd3; 23344: data <= 'd3; 23345: data <= 'd3; 23346: data <= 'd3; 23347: data <= 'd1; 23348: data <= 'd1; 23349: data <= 'd4; 23350: data <= 'd2; 23351: data <= 'd0; 23352: data <= 'd0; 23353: data <= 'd0; 23354: data <= 'd0; 23355: data <= 'd0; 23356: data <= 'd0; 23357: data <= 'd0; 23358: data <= 'd0; 23359: data <= 'd0; 23360: data <= 'd0; 23361: data <= 'd0; 23362: data <= 'd0; 23363: data <= 'd0; 23364: data <= 'd0; 23365: data <= 'd0; 23366: data <= 'd0; 23367: data <= 'd2; 23368: data <= 'd10; 23369: data <= 'd10; 23370: data <= 'd2; 23371: data <= 'd1; 23372: data <= 'd1; 23373: data <= 'd3; 23374: data <= 'd3; 23375: data <= 'd3; 23376: data <= 'd3; 23377: data <= 'd3; 23378: data <= 'd1; 23379: data <= 'd1; 23380: data <= 'd2; 23381: data <= 'd10; 23382: data <= 'd10; 23383: data <= 'd2; 23384: data <= 'd0; 23385: data <= 'd0; 23386: data <= 'd0; 23387: data <= 'd0; 23388: data <= 'd0; 23389: data <= 'd0; 23390: data <= 'd0; 23391: data <= 'd0; 23392: data <= 'd0; 23393: data <= 'd0; 23394: data <= 'd0; 23395: data <= 'd0; 23396: data <= 'd0; 23397: data <= 'd0; 23398: data <= 'd0; 23399: data <= 'd2; 23400: data <= 'd10; 23401: data <= 'd10; 23402: data <= 'd2; 23403: data <= 'd2; 23404: data <= 'd2; 23405: data <= 'd2; 23406: data <= 'd5; 23407: data <= 'd5; 23408: data <= 'd5; 23409: data <= 'd2; 23410: data <= 'd2; 23411: data <= 'd2; 23412: data <= 'd2; 23413: data <= 'd10; 23414: data <= 'd10; 23415: data <= 'd2; 23416: data <= 'd0; 23417: data <= 'd0; 23418: data <= 'd0; 23419: data <= 'd0; 23420: data <= 'd0; 23421: data <= 'd0; 23422: data <= 'd0; 23423: data <= 'd0; 23424: data <= 'd0; 23425: data <= 'd0; 23426: data <= 'd0; 23427: data <= 'd0; 23428: data <= 'd0; 23429: data <= 'd0; 23430: data <= 'd0; 23431: data <= 'd0; 23432: data <= 'd2; 23433: data <= 'd2; 23434: data <= 'd2; 23435: data <= 'd1; 23436: data <= 'd1; 23437: data <= 'd3; 23438: data <= 'd3; 23439: data <= 'd3; 23440: data <= 'd3; 23441: data <= 'd3; 23442: data <= 'd1; 23443: data <= 'd1; 23444: data <= 'd2; 23445: data <= 'd2; 23446: data <= 'd2; 23447: data <= 'd0; 23448: data <= 'd0; 23449: data <= 'd0; 23450: data <= 'd0; 23451: data <= 'd0; 23452: data <= 'd0; 23453: data <= 'd0; 23454: data <= 'd0; 23455: data <= 'd0; 23456: data <= 'd0; 23457: data <= 'd0; 23458: data <= 'd0; 23459: data <= 'd0; 23460: data <= 'd0; 23461: data <= 'd0; 23462: data <= 'd0; 23463: data <= 'd0; 23464: data <= 'd0; 23465: data <= 'd0; 23466: data <= 'd2; 23467: data <= 'd7; 23468: data <= 'd7; 23469: data <= 'd4; 23470: data <= 'd2; 23471: data <= 'd2; 23472: data <= 'd2; 23473: data <= 'd4; 23474: data <= 'd7; 23475: data <= 'd7; 23476: data <= 'd2; 23477: data <= 'd0; 23478: data <= 'd0; 23479: data <= 'd0; 23480: data <= 'd0; 23481: data <= 'd0; 23482: data <= 'd0; 23483: data <= 'd0; 23484: data <= 'd0; 23485: data <= 'd0; 23486: data <= 'd0; 23487: data <= 'd0; 23488: data <= 'd0; 23489: data <= 'd0; 23490: data <= 'd0; 23491: data <= 'd0; 23492: data <= 'd0; 23493: data <= 'd0; 23494: data <= 'd0; 23495: data <= 'd0; 23496: data <= 'd0; 23497: data <= 'd0; 23498: data <= 'd2; 23499: data <= 'd7; 23500: data <= 'd4; 23501: data <= 'd2; 23502: data <= 'd0; 23503: data <= 'd0; 23504: data <= 'd0; 23505: data <= 'd2; 23506: data <= 'd4; 23507: data <= 'd7; 23508: data <= 'd2; 23509: data <= 'd0; 23510: data <= 'd0; 23511: data <= 'd0; 23512: data <= 'd0; 23513: data <= 'd0; 23514: data <= 'd0; 23515: data <= 'd0; 23516: data <= 'd0; 23517: data <= 'd0; 23518: data <= 'd0; 23519: data <= 'd0; 23520: data <= 'd0; 23521: data <= 'd0; 23522: data <= 'd0; 23523: data <= 'd0; 23524: data <= 'd0; 23525: data <= 'd0; 23526: data <= 'd0; 23527: data <= 'd0; 23528: data <= 'd0; 23529: data <= 'd0; 23530: data <= 'd2; 23531: data <= 'd2; 23532: data <= 'd2; 23533: data <= 'd0; 23534: data <= 'd0; 23535: data <= 'd0; 23536: data <= 'd0; 23537: data <= 'd0; 23538: data <= 'd2; 23539: data <= 'd2; 23540: data <= 'd2; 23541: data <= 'd0; 23542: data <= 'd0; 23543: data <= 'd0; 23544: data <= 'd0; 23545: data <= 'd0; 23546: data <= 'd0; 23547: data <= 'd0; 23548: data <= 'd0; 23549: data <= 'd0; 23550: data <= 'd0; 23551: data <= 'd0;         
        endcase
    end
assign dout = data;

endmodule