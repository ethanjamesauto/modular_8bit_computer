module instruction_decoder(
);