// ROMs Using Block RAM Resources.
// File: rams_sp_rom_1.v
//
module ground_tex_rom(clk, en, addr, dout);
input clk;
input en;
input [7:0] addr;
output [2:0] dout;

logic [2:0] data;

always_ff @(posedge clk) begin
    if (en)
        case(addr)
            0: data <= 3'd4;1: data <= 3'd4;2: data <= 3'd4;3: data <= 3'd1;4: data <= 3'd4;5: data <= 3'd4;6: data <= 3'd2;7: data <= 3'd4;8: data <= 3'd1;9: data <= 3'd2;10: data <= 3'd4;11: data <= 3'd4;12: data <= 3'd4;13: data <= 3'd1;14: data <= 3'd2;15: data <= 3'd1;16: data <= 3'd1;17: data <= 3'd1;18: data <= 3'd1;19: data <= 3'd2;20: data <= 3'd1;21: data <= 3'd1;22: data <= 3'd2;23: data <= 3'd1;24: data <= 3'd2;25: data <= 3'd3;26: data <= 3'd1;27: data <= 3'd1;28: data <= 3'd1;29: data <= 3'd1;30: data <= 3'd2;31: data <= 3'd1;32: data <= 3'd1;33: data <= 3'd2;34: data <= 3'd3;35: data <= 3'd3;36: data <= 3'd2;37: data <= 3'd1;38: data <= 3'd3;39: data <= 3'd3;40: data <= 3'd7;41: data <= 3'd3;42: data <= 3'd2;43: data <= 3'd1;44: data <= 3'd2;45: data <= 3'd3;46: data <= 3'd3;47: data <= 3'd2;48: data <= 3'd3;49: data <= 3'd3;50: data <= 3'd3;51: data <= 3'd5;52: data <= 3'd5;53: data <= 3'd2;54: data <= 3'd3;55: data <= 3'd6;56: data <= 3'd6;57: data <= 3'd6;58: data <= 3'd3;59: data <= 3'd3;60: data <= 3'd6;61: data <= 3'd6;62: data <= 3'd6;63: data <= 3'd3;64: data <= 3'd5;65: data <= 3'd6;66: data <= 3'd6;67: data <= 3'd5;68: data <= 3'd3;69: data <= 3'd3;70: data <= 3'd5;71: data <= 3'd6;72: data <= 3'd6;73: data <= 3'd5;74: data <= 3'd3;75: data <= 3'd3;76: data <= 3'd5;77: data <= 3'd6;78: data <= 3'd6;79: data <= 3'd5;80: data <= 3'd0;81: data <= 3'd5;82: data <= 3'd5;83: data <= 3'd3;84: data <= 3'd0;85: data <= 3'd5;86: data <= 3'd5;87: data <= 3'd3;88: data <= 3'd5;89: data <= 3'd3;90: data <= 3'd5;91: data <= 3'd5;92: data <= 3'd3;93: data <= 3'd5;94: data <= 3'd5;95: data <= 3'd0;96: data <= 3'd0;97: data <= 3'd3;98: data <= 3'd3;99: data <= 3'd3;100: data <= 3'd0;101: data <= 3'd3;102: data <= 3'd3;103: data <= 3'd0;104: data <= 3'd3;105: data <= 3'd0;106: data <= 3'd5;107: data <= 3'd5;108: data <= 3'd0;109: data <= 3'd3;110: data <= 3'd3;111: data <= 3'd0;112: data <= 3'd3;113: data <= 3'd0;114: data <= 3'd3;115: data <= 3'd3;116: data <= 3'd0;117: data <= 3'd0;118: data <= 3'd0;119: data <= 3'd0;120: data <= 3'd0;121: data <= 3'd0;122: data <= 3'd3;123: data <= 3'd3;124: data <= 3'd0;125: data <= 3'd3;126: data <= 3'd0;127: data <= 3'd3;128: data <= 3'd3;129: data <= 3'd0;130: data <= 3'd0;131: data <= 3'd0;132: data <= 3'd0;133: data <= 3'd0;134: data <= 3'd0;135: data <= 3'd3;136: data <= 3'd0;137: data <= 3'd0;138: data <= 3'd0;139: data <= 3'd0;140: data <= 3'd0;141: data <= 3'd0;142: data <= 3'd0;143: data <= 3'd3;144: data <= 3'd0;145: data <= 3'd0;146: data <= 3'd0;147: data <= 3'd0;148: data <= 3'd0;149: data <= 3'd0;150: data <= 3'd0;151: data <= 3'd0;152: data <= 3'd0;153: data <= 3'd0;154: data <= 3'd0;155: data <= 3'd0;156: data <= 3'd0;157: data <= 3'd0;158: data <= 3'd0;159: data <= 3'd0;160: data <= 3'd0;161: data <= 3'd0;162: data <= 3'd0;163: data <= 3'd0;164: data <= 3'd0;165: data <= 3'd0;166: data <= 3'd0;167: data <= 3'd0;168: data <= 3'd0;169: data <= 3'd0;170: data <= 3'd0;171: data <= 3'd0;172: data <= 3'd0;173: data <= 3'd0;174: data <= 3'd0;175: data <= 3'd0;176: data <= 3'd0;177: data <= 3'd0;178: data <= 3'd0;179: data <= 3'd0;180: data <= 3'd0;181: data <= 3'd0;182: data <= 3'd0;183: data <= 3'd0;184: data <= 3'd0;185: data <= 3'd0;186: data <= 3'd0;187: data <= 3'd0;188: data <= 3'd0;189: data <= 3'd0;190: data <= 3'd0;191: data <= 3'd0;192: data <= 3'd0;193: data <= 3'd0;194: data <= 3'd0;195: data <= 3'd0;196: data <= 3'd0;197: data <= 3'd0;198: data <= 3'd0;199: data <= 3'd0;200: data <= 3'd0;201: data <= 3'd0;202: data <= 3'd0;203: data <= 3'd0;204: data <= 3'd0;205: data <= 3'd0;206: data <= 3'd0;207: data <= 3'd0;208: data <= 3'd0;209: data <= 3'd0;210: data <= 3'd0;211: data <= 3'd0;212: data <= 3'd0;213: data <= 3'd0;214: data <= 3'd0;215: data <= 3'd0;216: data <= 3'd0;217: data <= 3'd0;218: data <= 3'd0;219: data <= 3'd0;220: data <= 3'd0;221: data <= 3'd0;222: data <= 3'd0;223: data <= 3'd0;224: data <= 3'd0;225: data <= 3'd0;226: data <= 3'd0;227: data <= 3'd0;228: data <= 3'd0;229: data <= 3'd0;230: data <= 3'd0;231: data <= 3'd0;232: data <= 3'd0;233: data <= 3'd0;234: data <= 3'd0;235: data <= 3'd0;236: data <= 3'd0;237: data <= 3'd0;238: data <= 3'd0;239: data <= 3'd0;240: data <= 3'd0;241: data <= 3'd0;242: data <= 3'd0;243: data <= 3'd0;244: data <= 3'd0;245: data <= 3'd0;246: data <= 3'd0;247: data <= 3'd0;248: data <= 3'd0;249: data <= 3'd0;250: data <= 3'd0;251: data <= 3'd0;252: data <= 3'd0;253: data <= 3'd0;254: data <= 3'd0;255: data <= 3'd0;
        endcase
    end
assign dout = data;

endmodule