// This module models the computer as a whole
// and as such has no IOs. However, future IOs may be
// added for simulating user IO.
`timescale 1us/1us

module top;


// Below are any wires from card external
// IO for debugging purposes
// (nothing here right now)


// The main bus wires (32+8=40 wires total)
// On the bus connector, all buses have LSBs closer to the power pins and MSBs farther away
wire VCC_5V;
wire GND;
wire clk;			      // generated by motherboard clock generator
wire rst_n;			    // probably a button on the motherboard
wire VCC_3V3;
wire we_n;			      // active LOW
wire oe_n;			      // active LOW
wire int_n;			    // pulled up by motherboard; driven down by any peripheral (could be used for interrupts)
wire [7:0] data;
wire [15:0] addr;	  // 64k address space is suppored by default. More address bits may be added later
wire [7:0] aux_bus;

// Below are where test cards are instantiated
simple_card simple_card0(
	.VCC(VCC),
	.GND(GND),
	.clk(clk),
	.rst_n(rst_n),
	.we_n(we_n),
	.oe_n(oe_n),
	.data(data),
	.addr(addr),
	.int_n(int_n)
);

cpu_card cpu_card0(
	.VCC(VCC),
	.GND(GND),
	.clk(clk),
	.rst_n(rst_n),
	.we_n(we_n),
	.oe_n(oe_n),
	.data(data),
	.addr(addr),
	.int_n(int_n)
);

alu_card alu_card0(
	.VCC(VCC),
	.GND(GND),
	.clk(clk),
	.rst_n(rst_n),
	.we_n(we_n),
	.oe_n(oe_n),
	.data(data),
	.addr(addr),
	.int_n(int_n)
);

/*
module shift_card(
    input wire VCC,
    input wire GND,
    input wire clk,				// generated by motherboard clock generator
    input wire rst_n,			// probably a button on the motherboard
    input reg we_n,			    // active low
    input reg oe_n,			    // active low
    inout wire [7:0] data,
    input wire [15:0] addr,	    // 64k address space is suppored by default. More address bits may be added later
    output wire int_n,			// pulled up by motherboard; driven down by any peripheral (could be used for interrupts)
    output wire [7:0] aux_bus,
    output reg [7:0] TO_BUFFER_DATA,
    output wire TO_BUFFER_OE_N,
    output wire TO_AUX_BUS
);
*/

wire TO_BUFFER_DATA;
wire TO_BUFFER_DATA_OE_N;
wire TO_AUX_BUS;

shift_card shift_card0(
	.VCC(VCC),
	.GND(GND),
	.clk(clk),
	.rst_n(rst_n),
	.we_n(we_n),
	.oe_n(oe_n),
	.data(data),
	.addr(addr),
	.int_n(int_n),
	.aux_bus(aux_bus),
	.TO_BUFFER_DATA(TO_BUFFER_DATA),
	.TO_BUFFER_OE_N(TO_BUFFER_DATA_OE_N),
	.TO_AUX_BUS(TO_AUX_BUS)
);

// Below is motherboard logic (most of it is simulated and non-synthesizable)
assign VCC = 1'b1;
assign GND = 1'b0;

pullup(int_n);

reg clk_gen, rst_n_gen;
assign clk = clk_gen;
assign rst_n = rst_n_gen;

// clock
initial begin
	clk_gen = 1'b0;
	forever #1 clk_gen = ~clk_gen;
end

// reset
initial begin
	rst_n_gen = 1'b1;
	#2 rst_n_gen = 1'b0;
	#2 rst_n_gen = 1'b1;
end

endmodule